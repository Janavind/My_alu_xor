magic
tech sky130A
magscale 1 2
timestamp 1647379109
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 750 2128 178848 118992
<< metal2 >>
rect 754 119200 810 120000
rect 2226 119200 2282 120000
rect 3698 119200 3754 120000
rect 5262 119200 5318 120000
rect 6734 119200 6790 120000
rect 8298 119200 8354 120000
rect 9770 119200 9826 120000
rect 11334 119200 11390 120000
rect 12806 119200 12862 120000
rect 14370 119200 14426 120000
rect 15842 119200 15898 120000
rect 17314 119200 17370 120000
rect 18878 119200 18934 120000
rect 20350 119200 20406 120000
rect 21914 119200 21970 120000
rect 23386 119200 23442 120000
rect 24950 119200 25006 120000
rect 26422 119200 26478 120000
rect 27986 119200 28042 120000
rect 29458 119200 29514 120000
rect 30930 119200 30986 120000
rect 32494 119200 32550 120000
rect 33966 119200 34022 120000
rect 35530 119200 35586 120000
rect 37002 119200 37058 120000
rect 38566 119200 38622 120000
rect 40038 119200 40094 120000
rect 41602 119200 41658 120000
rect 43074 119200 43130 120000
rect 44546 119200 44602 120000
rect 46110 119200 46166 120000
rect 47582 119200 47638 120000
rect 49146 119200 49202 120000
rect 50618 119200 50674 120000
rect 52182 119200 52238 120000
rect 53654 119200 53710 120000
rect 55218 119200 55274 120000
rect 56690 119200 56746 120000
rect 58162 119200 58218 120000
rect 59726 119200 59782 120000
rect 61198 119200 61254 120000
rect 62762 119200 62818 120000
rect 64234 119200 64290 120000
rect 65798 119200 65854 120000
rect 67270 119200 67326 120000
rect 68834 119200 68890 120000
rect 70306 119200 70362 120000
rect 71778 119200 71834 120000
rect 73342 119200 73398 120000
rect 74814 119200 74870 120000
rect 76378 119200 76434 120000
rect 77850 119200 77906 120000
rect 79414 119200 79470 120000
rect 80886 119200 80942 120000
rect 82450 119200 82506 120000
rect 83922 119200 83978 120000
rect 85394 119200 85450 120000
rect 86958 119200 87014 120000
rect 88430 119200 88486 120000
rect 89994 119200 90050 120000
rect 91466 119200 91522 120000
rect 93030 119200 93086 120000
rect 94502 119200 94558 120000
rect 96066 119200 96122 120000
rect 97538 119200 97594 120000
rect 99010 119200 99066 120000
rect 100574 119200 100630 120000
rect 102046 119200 102102 120000
rect 103610 119200 103666 120000
rect 105082 119200 105138 120000
rect 106646 119200 106702 120000
rect 108118 119200 108174 120000
rect 109682 119200 109738 120000
rect 111154 119200 111210 120000
rect 112626 119200 112682 120000
rect 114190 119200 114246 120000
rect 115662 119200 115718 120000
rect 117226 119200 117282 120000
rect 118698 119200 118754 120000
rect 120262 119200 120318 120000
rect 121734 119200 121790 120000
rect 123298 119200 123354 120000
rect 124770 119200 124826 120000
rect 126242 119200 126298 120000
rect 127806 119200 127862 120000
rect 129278 119200 129334 120000
rect 130842 119200 130898 120000
rect 132314 119200 132370 120000
rect 133878 119200 133934 120000
rect 135350 119200 135406 120000
rect 136914 119200 136970 120000
rect 138386 119200 138442 120000
rect 139858 119200 139914 120000
rect 141422 119200 141478 120000
rect 142894 119200 142950 120000
rect 144458 119200 144514 120000
rect 145930 119200 145986 120000
rect 147494 119200 147550 120000
rect 148966 119200 149022 120000
rect 150530 119200 150586 120000
rect 152002 119200 152058 120000
rect 153474 119200 153530 120000
rect 155038 119200 155094 120000
rect 156510 119200 156566 120000
rect 158074 119200 158130 120000
rect 159546 119200 159602 120000
rect 161110 119200 161166 120000
rect 162582 119200 162638 120000
rect 164146 119200 164202 120000
rect 165618 119200 165674 120000
rect 167090 119200 167146 120000
rect 168654 119200 168710 120000
rect 170126 119200 170182 120000
rect 171690 119200 171746 120000
rect 173162 119200 173218 120000
rect 174726 119200 174782 120000
rect 176198 119200 176254 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31758 0 31814 800
rect 32126 0 32182 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44638 0 44694 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45742 0 45798 800
rect 46018 0 46074 800
rect 46386 0 46442 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47858 0 47914 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53194 0 53250 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56414 0 56470 800
rect 56782 0 56838 800
rect 57150 0 57206 800
rect 57426 0 57482 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65706 0 65762 800
rect 65982 0 66038 800
rect 66350 0 66406 800
rect 66718 0 66774 800
rect 67086 0 67142 800
rect 67454 0 67510 800
rect 67822 0 67878 800
rect 68190 0 68246 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69570 0 69626 800
rect 69938 0 69994 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80242 0 80298 800
rect 80610 0 80666 800
rect 80978 0 81034 800
rect 81346 0 81402 800
rect 81714 0 81770 800
rect 82082 0 82138 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83094 0 83150 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84198 0 84254 800
rect 84566 0 84622 800
rect 84934 0 84990 800
rect 85302 0 85358 800
rect 85670 0 85726 800
rect 85946 0 86002 800
rect 86314 0 86370 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87418 0 87474 800
rect 87786 0 87842 800
rect 88154 0 88210 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91650 0 91706 800
rect 92018 0 92074 800
rect 92386 0 92442 800
rect 92754 0 92810 800
rect 93122 0 93178 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94226 0 94282 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95238 0 95294 800
rect 95606 0 95662 800
rect 95974 0 96030 800
rect 96342 0 96398 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97354 0 97410 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98458 0 98514 800
rect 98826 0 98882 800
rect 99194 0 99250 800
rect 99562 0 99618 800
rect 99930 0 99986 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 105910 0 105966 800
rect 106278 0 106334 800
rect 106646 0 106702 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107750 0 107806 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109498 0 109554 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111338 0 111394 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112718 0 112774 800
rect 113086 0 113142 800
rect 113454 0 113510 800
rect 113822 0 113878 800
rect 114190 0 114246 800
rect 114466 0 114522 800
rect 114834 0 114890 800
rect 115202 0 115258 800
rect 115570 0 115626 800
rect 115938 0 115994 800
rect 116306 0 116362 800
rect 116674 0 116730 800
rect 117042 0 117098 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 118054 0 118110 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124126 0 124182 800
rect 124494 0 124550 800
rect 124862 0 124918 800
rect 125230 0 125286 800
rect 125598 0 125654 800
rect 125874 0 125930 800
rect 126242 0 126298 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127346 0 127402 800
rect 127714 0 127770 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130566 0 130622 800
rect 130934 0 130990 800
rect 131302 0 131358 800
rect 131578 0 131634 800
rect 131946 0 132002 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134430 0 134486 800
rect 134798 0 134854 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 137006 0 137062 800
rect 137282 0 137338 800
rect 137650 0 137706 800
rect 138018 0 138074 800
rect 138386 0 138442 800
rect 138754 0 138810 800
rect 139122 0 139178 800
rect 139490 0 139546 800
rect 139858 0 139914 800
rect 140134 0 140190 800
rect 140502 0 140558 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141606 0 141662 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143722 0 143778 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145838 0 145894 800
rect 146206 0 146262 800
rect 146574 0 146630 800
rect 146942 0 146998 800
rect 147310 0 147366 800
rect 147678 0 147734 800
rect 148046 0 148102 800
rect 148414 0 148470 800
rect 148690 0 148746 800
rect 149058 0 149114 800
rect 149426 0 149482 800
rect 149794 0 149850 800
rect 150162 0 150218 800
rect 150530 0 150586 800
rect 150898 0 150954 800
rect 151266 0 151322 800
rect 151542 0 151598 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152646 0 152702 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153750 0 153806 800
rect 154118 0 154174 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157246 0 157302 800
rect 157614 0 157670 800
rect 157982 0 158038 800
rect 158350 0 158406 800
rect 158718 0 158774 800
rect 159086 0 159142 800
rect 159454 0 159510 800
rect 159822 0 159878 800
rect 160098 0 160154 800
rect 160466 0 160522 800
rect 160834 0 160890 800
rect 161202 0 161258 800
rect 161570 0 161626 800
rect 161938 0 161994 800
rect 162306 0 162362 800
rect 162674 0 162730 800
rect 162950 0 163006 800
rect 163318 0 163374 800
rect 163686 0 163742 800
rect 164054 0 164110 800
rect 164422 0 164478 800
rect 164790 0 164846 800
rect 165158 0 165214 800
rect 165526 0 165582 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 168010 0 168066 800
rect 168378 0 168434 800
rect 168654 0 168710 800
rect 169022 0 169078 800
rect 169390 0 169446 800
rect 169758 0 169814 800
rect 170126 0 170182 800
rect 170494 0 170550 800
rect 170862 0 170918 800
rect 171230 0 171286 800
rect 171506 0 171562 800
rect 171874 0 171930 800
rect 172242 0 172298 800
rect 172610 0 172666 800
rect 172978 0 173034 800
rect 173346 0 173402 800
rect 173714 0 173770 800
rect 174082 0 174138 800
rect 174358 0 174414 800
rect 174726 0 174782 800
rect 175094 0 175150 800
rect 175462 0 175518 800
rect 175830 0 175886 800
rect 176198 0 176254 800
rect 176566 0 176622 800
rect 176934 0 176990 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 866 119144 2170 119354
rect 2338 119144 3642 119354
rect 3810 119144 5206 119354
rect 5374 119144 6678 119354
rect 6846 119144 8242 119354
rect 8410 119144 9714 119354
rect 9882 119144 11278 119354
rect 11446 119144 12750 119354
rect 12918 119144 14314 119354
rect 14482 119144 15786 119354
rect 15954 119144 17258 119354
rect 17426 119144 18822 119354
rect 18990 119144 20294 119354
rect 20462 119144 21858 119354
rect 22026 119144 23330 119354
rect 23498 119144 24894 119354
rect 25062 119144 26366 119354
rect 26534 119144 27930 119354
rect 28098 119144 29402 119354
rect 29570 119144 30874 119354
rect 31042 119144 32438 119354
rect 32606 119144 33910 119354
rect 34078 119144 35474 119354
rect 35642 119144 36946 119354
rect 37114 119144 38510 119354
rect 38678 119144 39982 119354
rect 40150 119144 41546 119354
rect 41714 119144 43018 119354
rect 43186 119144 44490 119354
rect 44658 119144 46054 119354
rect 46222 119144 47526 119354
rect 47694 119144 49090 119354
rect 49258 119144 50562 119354
rect 50730 119144 52126 119354
rect 52294 119144 53598 119354
rect 53766 119144 55162 119354
rect 55330 119144 56634 119354
rect 56802 119144 58106 119354
rect 58274 119144 59670 119354
rect 59838 119144 61142 119354
rect 61310 119144 62706 119354
rect 62874 119144 64178 119354
rect 64346 119144 65742 119354
rect 65910 119144 67214 119354
rect 67382 119144 68778 119354
rect 68946 119144 70250 119354
rect 70418 119144 71722 119354
rect 71890 119144 73286 119354
rect 73454 119144 74758 119354
rect 74926 119144 76322 119354
rect 76490 119144 77794 119354
rect 77962 119144 79358 119354
rect 79526 119144 80830 119354
rect 80998 119144 82394 119354
rect 82562 119144 83866 119354
rect 84034 119144 85338 119354
rect 85506 119144 86902 119354
rect 87070 119144 88374 119354
rect 88542 119144 89938 119354
rect 90106 119144 91410 119354
rect 91578 119144 92974 119354
rect 93142 119144 94446 119354
rect 94614 119144 96010 119354
rect 96178 119144 97482 119354
rect 97650 119144 98954 119354
rect 99122 119144 100518 119354
rect 100686 119144 101990 119354
rect 102158 119144 103554 119354
rect 103722 119144 105026 119354
rect 105194 119144 106590 119354
rect 106758 119144 108062 119354
rect 108230 119144 109626 119354
rect 109794 119144 111098 119354
rect 111266 119144 112570 119354
rect 112738 119144 114134 119354
rect 114302 119144 115606 119354
rect 115774 119144 117170 119354
rect 117338 119144 118642 119354
rect 118810 119144 120206 119354
rect 120374 119144 121678 119354
rect 121846 119144 123242 119354
rect 123410 119144 124714 119354
rect 124882 119144 126186 119354
rect 126354 119144 127750 119354
rect 127918 119144 129222 119354
rect 129390 119144 130786 119354
rect 130954 119144 132258 119354
rect 132426 119144 133822 119354
rect 133990 119144 135294 119354
rect 135462 119144 136858 119354
rect 137026 119144 138330 119354
rect 138498 119144 139802 119354
rect 139970 119144 141366 119354
rect 141534 119144 142838 119354
rect 143006 119144 144402 119354
rect 144570 119144 145874 119354
rect 146042 119144 147438 119354
rect 147606 119144 148910 119354
rect 149078 119144 150474 119354
rect 150642 119144 151946 119354
rect 152114 119144 153418 119354
rect 153586 119144 154982 119354
rect 155150 119144 156454 119354
rect 156622 119144 158018 119354
rect 158186 119144 159490 119354
rect 159658 119144 161054 119354
rect 161222 119144 162526 119354
rect 162694 119144 164090 119354
rect 164258 119144 165562 119354
rect 165730 119144 167034 119354
rect 167202 119144 168598 119354
rect 168766 119144 170070 119354
rect 170238 119144 171634 119354
rect 171802 119144 173106 119354
rect 173274 119144 174670 119354
rect 174838 119144 175516 119354
rect 756 856 175516 119144
rect 866 800 1066 856
rect 1234 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3182 856
rect 3350 800 3550 856
rect 3718 800 3918 856
rect 4086 800 4286 856
rect 4454 800 4654 856
rect 4822 800 5022 856
rect 5190 800 5390 856
rect 5558 800 5758 856
rect 5926 800 6034 856
rect 6202 800 6402 856
rect 6570 800 6770 856
rect 6938 800 7138 856
rect 7306 800 7506 856
rect 7674 800 7874 856
rect 8042 800 8242 856
rect 8410 800 8610 856
rect 8778 800 8886 856
rect 9054 800 9254 856
rect 9422 800 9622 856
rect 9790 800 9990 856
rect 10158 800 10358 856
rect 10526 800 10726 856
rect 10894 800 11094 856
rect 11262 800 11462 856
rect 11630 800 11738 856
rect 11906 800 12106 856
rect 12274 800 12474 856
rect 12642 800 12842 856
rect 13010 800 13210 856
rect 13378 800 13578 856
rect 13746 800 13946 856
rect 14114 800 14314 856
rect 14482 800 14590 856
rect 14758 800 14958 856
rect 15126 800 15326 856
rect 15494 800 15694 856
rect 15862 800 16062 856
rect 16230 800 16430 856
rect 16598 800 16798 856
rect 16966 800 17166 856
rect 17334 800 17442 856
rect 17610 800 17810 856
rect 17978 800 18178 856
rect 18346 800 18546 856
rect 18714 800 18914 856
rect 19082 800 19282 856
rect 19450 800 19650 856
rect 19818 800 20018 856
rect 20186 800 20294 856
rect 20462 800 20662 856
rect 20830 800 21030 856
rect 21198 800 21398 856
rect 21566 800 21766 856
rect 21934 800 22134 856
rect 22302 800 22502 856
rect 22670 800 22870 856
rect 23038 800 23146 856
rect 23314 800 23514 856
rect 23682 800 23882 856
rect 24050 800 24250 856
rect 24418 800 24618 856
rect 24786 800 24986 856
rect 25154 800 25354 856
rect 25522 800 25722 856
rect 25890 800 25998 856
rect 26166 800 26366 856
rect 26534 800 26734 856
rect 26902 800 27102 856
rect 27270 800 27470 856
rect 27638 800 27838 856
rect 28006 800 28206 856
rect 28374 800 28574 856
rect 28742 800 28850 856
rect 29018 800 29218 856
rect 29386 800 29586 856
rect 29754 800 29954 856
rect 30122 800 30322 856
rect 30490 800 30690 856
rect 30858 800 31058 856
rect 31226 800 31426 856
rect 31594 800 31702 856
rect 31870 800 32070 856
rect 32238 800 32438 856
rect 32606 800 32806 856
rect 32974 800 33174 856
rect 33342 800 33542 856
rect 33710 800 33910 856
rect 34078 800 34278 856
rect 34446 800 34554 856
rect 34722 800 34922 856
rect 35090 800 35290 856
rect 35458 800 35658 856
rect 35826 800 36026 856
rect 36194 800 36394 856
rect 36562 800 36762 856
rect 36930 800 37130 856
rect 37298 800 37406 856
rect 37574 800 37774 856
rect 37942 800 38142 856
rect 38310 800 38510 856
rect 38678 800 38878 856
rect 39046 800 39246 856
rect 39414 800 39614 856
rect 39782 800 39982 856
rect 40150 800 40258 856
rect 40426 800 40626 856
rect 40794 800 40994 856
rect 41162 800 41362 856
rect 41530 800 41730 856
rect 41898 800 42098 856
rect 42266 800 42466 856
rect 42634 800 42834 856
rect 43002 800 43110 856
rect 43278 800 43478 856
rect 43646 800 43846 856
rect 44014 800 44214 856
rect 44382 800 44582 856
rect 44750 800 44950 856
rect 45118 800 45318 856
rect 45486 800 45686 856
rect 45854 800 45962 856
rect 46130 800 46330 856
rect 46498 800 46698 856
rect 46866 800 47066 856
rect 47234 800 47434 856
rect 47602 800 47802 856
rect 47970 800 48170 856
rect 48338 800 48538 856
rect 48706 800 48814 856
rect 48982 800 49182 856
rect 49350 800 49550 856
rect 49718 800 49918 856
rect 50086 800 50286 856
rect 50454 800 50654 856
rect 50822 800 51022 856
rect 51190 800 51390 856
rect 51558 800 51666 856
rect 51834 800 52034 856
rect 52202 800 52402 856
rect 52570 800 52770 856
rect 52938 800 53138 856
rect 53306 800 53506 856
rect 53674 800 53874 856
rect 54042 800 54242 856
rect 54410 800 54518 856
rect 54686 800 54886 856
rect 55054 800 55254 856
rect 55422 800 55622 856
rect 55790 800 55990 856
rect 56158 800 56358 856
rect 56526 800 56726 856
rect 56894 800 57094 856
rect 57262 800 57370 856
rect 57538 800 57738 856
rect 57906 800 58106 856
rect 58274 800 58474 856
rect 58642 800 58842 856
rect 59010 800 59210 856
rect 59378 800 59578 856
rect 59746 800 59946 856
rect 60114 800 60222 856
rect 60390 800 60590 856
rect 60758 800 60958 856
rect 61126 800 61326 856
rect 61494 800 61694 856
rect 61862 800 62062 856
rect 62230 800 62430 856
rect 62598 800 62798 856
rect 62966 800 63074 856
rect 63242 800 63442 856
rect 63610 800 63810 856
rect 63978 800 64178 856
rect 64346 800 64546 856
rect 64714 800 64914 856
rect 65082 800 65282 856
rect 65450 800 65650 856
rect 65818 800 65926 856
rect 66094 800 66294 856
rect 66462 800 66662 856
rect 66830 800 67030 856
rect 67198 800 67398 856
rect 67566 800 67766 856
rect 67934 800 68134 856
rect 68302 800 68502 856
rect 68670 800 68778 856
rect 68946 800 69146 856
rect 69314 800 69514 856
rect 69682 800 69882 856
rect 70050 800 70250 856
rect 70418 800 70618 856
rect 70786 800 70986 856
rect 71154 800 71354 856
rect 71522 800 71630 856
rect 71798 800 71998 856
rect 72166 800 72366 856
rect 72534 800 72734 856
rect 72902 800 73102 856
rect 73270 800 73470 856
rect 73638 800 73838 856
rect 74006 800 74206 856
rect 74374 800 74482 856
rect 74650 800 74850 856
rect 75018 800 75218 856
rect 75386 800 75586 856
rect 75754 800 75954 856
rect 76122 800 76322 856
rect 76490 800 76690 856
rect 76858 800 77058 856
rect 77226 800 77334 856
rect 77502 800 77702 856
rect 77870 800 78070 856
rect 78238 800 78438 856
rect 78606 800 78806 856
rect 78974 800 79174 856
rect 79342 800 79542 856
rect 79710 800 79910 856
rect 80078 800 80186 856
rect 80354 800 80554 856
rect 80722 800 80922 856
rect 81090 800 81290 856
rect 81458 800 81658 856
rect 81826 800 82026 856
rect 82194 800 82394 856
rect 82562 800 82762 856
rect 82930 800 83038 856
rect 83206 800 83406 856
rect 83574 800 83774 856
rect 83942 800 84142 856
rect 84310 800 84510 856
rect 84678 800 84878 856
rect 85046 800 85246 856
rect 85414 800 85614 856
rect 85782 800 85890 856
rect 86058 800 86258 856
rect 86426 800 86626 856
rect 86794 800 86994 856
rect 87162 800 87362 856
rect 87530 800 87730 856
rect 87898 800 88098 856
rect 88266 800 88466 856
rect 88634 800 88742 856
rect 88910 800 89110 856
rect 89278 800 89478 856
rect 89646 800 89846 856
rect 90014 800 90214 856
rect 90382 800 90582 856
rect 90750 800 90950 856
rect 91118 800 91318 856
rect 91486 800 91594 856
rect 91762 800 91962 856
rect 92130 800 92330 856
rect 92498 800 92698 856
rect 92866 800 93066 856
rect 93234 800 93434 856
rect 93602 800 93802 856
rect 93970 800 94170 856
rect 94338 800 94446 856
rect 94614 800 94814 856
rect 94982 800 95182 856
rect 95350 800 95550 856
rect 95718 800 95918 856
rect 96086 800 96286 856
rect 96454 800 96654 856
rect 96822 800 97022 856
rect 97190 800 97298 856
rect 97466 800 97666 856
rect 97834 800 98034 856
rect 98202 800 98402 856
rect 98570 800 98770 856
rect 98938 800 99138 856
rect 99306 800 99506 856
rect 99674 800 99874 856
rect 100042 800 100150 856
rect 100318 800 100518 856
rect 100686 800 100886 856
rect 101054 800 101254 856
rect 101422 800 101622 856
rect 101790 800 101990 856
rect 102158 800 102358 856
rect 102526 800 102726 856
rect 102894 800 103002 856
rect 103170 800 103370 856
rect 103538 800 103738 856
rect 103906 800 104106 856
rect 104274 800 104474 856
rect 104642 800 104842 856
rect 105010 800 105210 856
rect 105378 800 105578 856
rect 105746 800 105854 856
rect 106022 800 106222 856
rect 106390 800 106590 856
rect 106758 800 106958 856
rect 107126 800 107326 856
rect 107494 800 107694 856
rect 107862 800 108062 856
rect 108230 800 108430 856
rect 108598 800 108706 856
rect 108874 800 109074 856
rect 109242 800 109442 856
rect 109610 800 109810 856
rect 109978 800 110178 856
rect 110346 800 110546 856
rect 110714 800 110914 856
rect 111082 800 111282 856
rect 111450 800 111558 856
rect 111726 800 111926 856
rect 112094 800 112294 856
rect 112462 800 112662 856
rect 112830 800 113030 856
rect 113198 800 113398 856
rect 113566 800 113766 856
rect 113934 800 114134 856
rect 114302 800 114410 856
rect 114578 800 114778 856
rect 114946 800 115146 856
rect 115314 800 115514 856
rect 115682 800 115882 856
rect 116050 800 116250 856
rect 116418 800 116618 856
rect 116786 800 116986 856
rect 117154 800 117262 856
rect 117430 800 117630 856
rect 117798 800 117998 856
rect 118166 800 118366 856
rect 118534 800 118734 856
rect 118902 800 119102 856
rect 119270 800 119470 856
rect 119638 800 119838 856
rect 120006 800 120114 856
rect 120282 800 120482 856
rect 120650 800 120850 856
rect 121018 800 121218 856
rect 121386 800 121586 856
rect 121754 800 121954 856
rect 122122 800 122322 856
rect 122490 800 122690 856
rect 122858 800 122966 856
rect 123134 800 123334 856
rect 123502 800 123702 856
rect 123870 800 124070 856
rect 124238 800 124438 856
rect 124606 800 124806 856
rect 124974 800 125174 856
rect 125342 800 125542 856
rect 125710 800 125818 856
rect 125986 800 126186 856
rect 126354 800 126554 856
rect 126722 800 126922 856
rect 127090 800 127290 856
rect 127458 800 127658 856
rect 127826 800 128026 856
rect 128194 800 128394 856
rect 128562 800 128670 856
rect 128838 800 129038 856
rect 129206 800 129406 856
rect 129574 800 129774 856
rect 129942 800 130142 856
rect 130310 800 130510 856
rect 130678 800 130878 856
rect 131046 800 131246 856
rect 131414 800 131522 856
rect 131690 800 131890 856
rect 132058 800 132258 856
rect 132426 800 132626 856
rect 132794 800 132994 856
rect 133162 800 133362 856
rect 133530 800 133730 856
rect 133898 800 134098 856
rect 134266 800 134374 856
rect 134542 800 134742 856
rect 134910 800 135110 856
rect 135278 800 135478 856
rect 135646 800 135846 856
rect 136014 800 136214 856
rect 136382 800 136582 856
rect 136750 800 136950 856
rect 137118 800 137226 856
rect 137394 800 137594 856
rect 137762 800 137962 856
rect 138130 800 138330 856
rect 138498 800 138698 856
rect 138866 800 139066 856
rect 139234 800 139434 856
rect 139602 800 139802 856
rect 139970 800 140078 856
rect 140246 800 140446 856
rect 140614 800 140814 856
rect 140982 800 141182 856
rect 141350 800 141550 856
rect 141718 800 141918 856
rect 142086 800 142286 856
rect 142454 800 142654 856
rect 142822 800 142930 856
rect 143098 800 143298 856
rect 143466 800 143666 856
rect 143834 800 144034 856
rect 144202 800 144402 856
rect 144570 800 144770 856
rect 144938 800 145138 856
rect 145306 800 145506 856
rect 145674 800 145782 856
rect 145950 800 146150 856
rect 146318 800 146518 856
rect 146686 800 146886 856
rect 147054 800 147254 856
rect 147422 800 147622 856
rect 147790 800 147990 856
rect 148158 800 148358 856
rect 148526 800 148634 856
rect 148802 800 149002 856
rect 149170 800 149370 856
rect 149538 800 149738 856
rect 149906 800 150106 856
rect 150274 800 150474 856
rect 150642 800 150842 856
rect 151010 800 151210 856
rect 151378 800 151486 856
rect 151654 800 151854 856
rect 152022 800 152222 856
rect 152390 800 152590 856
rect 152758 800 152958 856
rect 153126 800 153326 856
rect 153494 800 153694 856
rect 153862 800 154062 856
rect 154230 800 154338 856
rect 154506 800 154706 856
rect 154874 800 155074 856
rect 155242 800 155442 856
rect 155610 800 155810 856
rect 155978 800 156178 856
rect 156346 800 156546 856
rect 156714 800 156914 856
rect 157082 800 157190 856
rect 157358 800 157558 856
rect 157726 800 157926 856
rect 158094 800 158294 856
rect 158462 800 158662 856
rect 158830 800 159030 856
rect 159198 800 159398 856
rect 159566 800 159766 856
rect 159934 800 160042 856
rect 160210 800 160410 856
rect 160578 800 160778 856
rect 160946 800 161146 856
rect 161314 800 161514 856
rect 161682 800 161882 856
rect 162050 800 162250 856
rect 162418 800 162618 856
rect 162786 800 162894 856
rect 163062 800 163262 856
rect 163430 800 163630 856
rect 163798 800 163998 856
rect 164166 800 164366 856
rect 164534 800 164734 856
rect 164902 800 165102 856
rect 165270 800 165470 856
rect 165638 800 165746 856
rect 165914 800 166114 856
rect 166282 800 166482 856
rect 166650 800 166850 856
rect 167018 800 167218 856
rect 167386 800 167586 856
rect 167754 800 167954 856
rect 168122 800 168322 856
rect 168490 800 168598 856
rect 168766 800 168966 856
rect 169134 800 169334 856
rect 169502 800 169702 856
rect 169870 800 170070 856
rect 170238 800 170438 856
rect 170606 800 170806 856
rect 170974 800 171174 856
rect 171342 800 171450 856
rect 171618 800 171818 856
rect 171986 800 172186 856
rect 172354 800 172554 856
rect 172722 800 172922 856
rect 173090 800 173290 856
rect 173458 800 173658 856
rect 173826 800 174026 856
rect 174194 800 174302 856
rect 174470 800 174670 856
rect 174838 800 175038 856
rect 175206 800 175406 856
<< metal3 >>
rect 0 109896 800 110016
rect 0 89904 800 90024
rect 0 69912 800 70032
rect 0 49920 800 50040
rect 0 29928 800 30048
rect 0 9936 800 10056
rect 179200 111392 180000 111512
rect 179200 94256 180000 94376
rect 179200 77120 180000 77240
rect 179200 59984 180000 60104
rect 179200 42848 180000 42968
rect 179200 25712 180000 25832
rect 179200 8576 180000 8696
<< obsm3 >>
rect 4208 2143 173488 118149
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 58203 117632 91389 118149
rect 58203 111691 65568 117632
rect 66048 111691 80928 117632
rect 81408 111691 91389 117632
<< labels >>
rlabel metal3 s 179200 8576 180000 8696 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 176198 119200 176254 120000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 179200 42848 180000 42968 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 179200 59984 180000 60104 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 177762 119200 177818 120000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 179200 77120 180000 77240 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 176566 0 176622 800 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 176934 0 176990 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 177210 0 177266 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 177578 0 177634 800 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 173162 119200 173218 120000 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 177946 0 178002 800 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 178314 0 178370 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 179200 94256 180000 94376 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 179200 111392 180000 111512 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 109896 800 110016 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 9936 800 10056 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 179200 25712 180000 25832 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 0 29928 800 30048 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 0 49920 800 50040 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 0 69912 800 70032 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal2 s 176198 0 176254 800 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 174726 119200 174782 120000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 0 89904 800 90024 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 30 nsew signal input
rlabel metal2 s 46110 119200 46166 120000 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 50618 119200 50674 120000 6 io_in[11]
port 32 nsew signal input
rlabel metal2 s 55218 119200 55274 120000 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 59726 119200 59782 120000 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 64234 119200 64290 120000 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 68834 119200 68890 120000 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 73342 119200 73398 120000 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 77850 119200 77906 120000 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 82450 119200 82506 120000 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 86958 119200 87014 120000 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 5262 119200 5318 120000 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 91466 119200 91522 120000 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 96066 119200 96122 120000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 100574 119200 100630 120000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 105082 119200 105138 120000 6 io_in[23]
port 45 nsew signal input
rlabel metal2 s 109682 119200 109738 120000 6 io_in[24]
port 46 nsew signal input
rlabel metal2 s 114190 119200 114246 120000 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 118698 119200 118754 120000 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 123298 119200 123354 120000 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 127806 119200 127862 120000 6 io_in[28]
port 50 nsew signal input
rlabel metal2 s 132314 119200 132370 120000 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 9770 119200 9826 120000 6 io_in[2]
port 52 nsew signal input
rlabel metal2 s 136914 119200 136970 120000 6 io_in[30]
port 53 nsew signal input
rlabel metal2 s 141422 119200 141478 120000 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 145930 119200 145986 120000 6 io_in[32]
port 55 nsew signal input
rlabel metal2 s 150530 119200 150586 120000 6 io_in[33]
port 56 nsew signal input
rlabel metal2 s 155038 119200 155094 120000 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 159546 119200 159602 120000 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 164146 119200 164202 120000 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 168654 119200 168710 120000 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 14370 119200 14426 120000 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 18878 119200 18934 120000 6 io_in[4]
port 62 nsew signal input
rlabel metal2 s 23386 119200 23442 120000 6 io_in[5]
port 63 nsew signal input
rlabel metal2 s 27986 119200 28042 120000 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 32494 119200 32550 120000 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 37002 119200 37058 120000 6 io_in[8]
port 66 nsew signal input
rlabel metal2 s 41602 119200 41658 120000 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 47582 119200 47638 120000 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 52182 119200 52238 120000 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 56690 119200 56746 120000 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 61198 119200 61254 120000 6 io_oeb[13]
port 72 nsew signal output
rlabel metal2 s 65798 119200 65854 120000 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 70306 119200 70362 120000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 74814 119200 74870 120000 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 79414 119200 79470 120000 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 83922 119200 83978 120000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 88430 119200 88486 120000 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 6734 119200 6790 120000 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 93030 119200 93086 120000 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 97538 119200 97594 120000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 102046 119200 102102 120000 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 106646 119200 106702 120000 6 io_oeb[23]
port 83 nsew signal output
rlabel metal2 s 111154 119200 111210 120000 6 io_oeb[24]
port 84 nsew signal output
rlabel metal2 s 115662 119200 115718 120000 6 io_oeb[25]
port 85 nsew signal output
rlabel metal2 s 120262 119200 120318 120000 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 124770 119200 124826 120000 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 129278 119200 129334 120000 6 io_oeb[28]
port 88 nsew signal output
rlabel metal2 s 133878 119200 133934 120000 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 11334 119200 11390 120000 6 io_oeb[2]
port 90 nsew signal output
rlabel metal2 s 138386 119200 138442 120000 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 142894 119200 142950 120000 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 147494 119200 147550 120000 6 io_oeb[32]
port 93 nsew signal output
rlabel metal2 s 152002 119200 152058 120000 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 156510 119200 156566 120000 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 161110 119200 161166 120000 6 io_oeb[35]
port 96 nsew signal output
rlabel metal2 s 165618 119200 165674 120000 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 170126 119200 170182 120000 6 io_oeb[37]
port 98 nsew signal output
rlabel metal2 s 15842 119200 15898 120000 6 io_oeb[3]
port 99 nsew signal output
rlabel metal2 s 20350 119200 20406 120000 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 24950 119200 25006 120000 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 29458 119200 29514 120000 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 33966 119200 34022 120000 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 38566 119200 38622 120000 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 43074 119200 43130 120000 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 3698 119200 3754 120000 6 io_out[0]
port 106 nsew signal output
rlabel metal2 s 49146 119200 49202 120000 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 53654 119200 53710 120000 6 io_out[11]
port 108 nsew signal output
rlabel metal2 s 58162 119200 58218 120000 6 io_out[12]
port 109 nsew signal output
rlabel metal2 s 62762 119200 62818 120000 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 67270 119200 67326 120000 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 71778 119200 71834 120000 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 76378 119200 76434 120000 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 80886 119200 80942 120000 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 85394 119200 85450 120000 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 89994 119200 90050 120000 6 io_out[19]
port 116 nsew signal output
rlabel metal2 s 8298 119200 8354 120000 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 94502 119200 94558 120000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 99010 119200 99066 120000 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 103610 119200 103666 120000 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 108118 119200 108174 120000 6 io_out[23]
port 121 nsew signal output
rlabel metal2 s 112626 119200 112682 120000 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 117226 119200 117282 120000 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 121734 119200 121790 120000 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 126242 119200 126298 120000 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 130842 119200 130898 120000 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 135350 119200 135406 120000 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 12806 119200 12862 120000 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 139858 119200 139914 120000 6 io_out[30]
port 129 nsew signal output
rlabel metal2 s 144458 119200 144514 120000 6 io_out[31]
port 130 nsew signal output
rlabel metal2 s 148966 119200 149022 120000 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 153474 119200 153530 120000 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 158074 119200 158130 120000 6 io_out[34]
port 133 nsew signal output
rlabel metal2 s 162582 119200 162638 120000 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 167090 119200 167146 120000 6 io_out[36]
port 135 nsew signal output
rlabel metal2 s 171690 119200 171746 120000 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 17314 119200 17370 120000 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 21914 119200 21970 120000 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 26422 119200 26478 120000 6 io_out[5]
port 139 nsew signal output
rlabel metal2 s 30930 119200 30986 120000 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 35530 119200 35586 120000 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 40038 119200 40094 120000 6 io_out[8]
port 142 nsew signal output
rlabel metal2 s 44546 119200 44602 120000 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 irq[0]
port 144 nsew signal output
rlabel metal2 s 175094 0 175150 800 6 irq[1]
port 145 nsew signal output
rlabel metal2 s 175462 0 175518 800 6 irq[2]
port 146 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 la_data_in[0]
port 147 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[100]
port 148 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_data_in[101]
port 149 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_data_in[102]
port 150 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_data_in[103]
port 151 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_data_in[104]
port 152 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_data_in[105]
port 153 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_data_in[106]
port 154 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[107]
port 155 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[108]
port 156 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_data_in[109]
port 157 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[10]
port 158 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[110]
port 159 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[111]
port 160 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 la_data_in[112]
port 161 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_data_in[113]
port 162 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_data_in[114]
port 163 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_data_in[115]
port 164 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_data_in[116]
port 165 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_data_in[117]
port 166 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_data_in[118]
port 167 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[119]
port 168 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[11]
port 169 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_data_in[120]
port 170 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_data_in[121]
port 171 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_data_in[122]
port 172 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 la_data_in[123]
port 173 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 la_data_in[124]
port 174 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_data_in[125]
port 175 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_data_in[126]
port 176 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_data_in[127]
port 177 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[12]
port 178 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_data_in[13]
port 179 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[14]
port 180 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[15]
port 181 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[16]
port 182 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[17]
port 183 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[18]
port 184 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[19]
port 185 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_data_in[1]
port 186 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[20]
port 187 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_data_in[21]
port 188 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[22]
port 189 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[23]
port 190 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[24]
port 191 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[25]
port 192 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[26]
port 193 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[27]
port 194 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[28]
port 195 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[29]
port 196 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[2]
port 197 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[30]
port 198 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[31]
port 199 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[32]
port 200 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[33]
port 201 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[34]
port 202 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[35]
port 203 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[36]
port 204 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[37]
port 205 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[38]
port 206 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[39]
port 207 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_data_in[3]
port 208 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[40]
port 209 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_data_in[41]
port 210 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[42]
port 211 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[43]
port 212 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[44]
port 213 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_data_in[45]
port 214 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[46]
port 215 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_data_in[47]
port 216 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[48]
port 217 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[49]
port 218 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_data_in[4]
port 219 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[50]
port 220 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[51]
port 221 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[52]
port 222 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[53]
port 223 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[54]
port 224 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[55]
port 225 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[56]
port 226 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[57]
port 227 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[58]
port 228 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[59]
port 229 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in[5]
port 230 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[60]
port 231 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[61]
port 232 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_data_in[62]
port 233 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[63]
port 234 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[64]
port 235 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[65]
port 236 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[66]
port 237 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[67]
port 238 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[68]
port 239 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_data_in[69]
port 240 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_data_in[6]
port 241 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[70]
port 242 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_data_in[71]
port 243 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[72]
port 244 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[73]
port 245 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[74]
port 246 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_data_in[75]
port 247 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[76]
port 248 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[77]
port 249 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_data_in[78]
port 250 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_data_in[79]
port 251 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[7]
port 252 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[80]
port 253 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_data_in[81]
port 254 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_data_in[82]
port 255 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_data_in[83]
port 256 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[84]
port 257 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_data_in[85]
port 258 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_data_in[86]
port 259 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_data_in[87]
port 260 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_data_in[88]
port 261 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_data_in[89]
port 262 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_data_in[8]
port 263 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 la_data_in[90]
port 264 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[91]
port 265 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[92]
port 266 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[93]
port 267 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_data_in[94]
port 268 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[95]
port 269 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_data_in[96]
port 270 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[97]
port 271 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_data_in[98]
port 272 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[99]
port 273 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[9]
port 274 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_data_out[0]
port 275 nsew signal output
rlabel metal2 s 145194 0 145250 800 6 la_data_out[100]
port 276 nsew signal output
rlabel metal2 s 146206 0 146262 800 6 la_data_out[101]
port 277 nsew signal output
rlabel metal2 s 147310 0 147366 800 6 la_data_out[102]
port 278 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 la_data_out[103]
port 279 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 la_data_out[104]
port 280 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[105]
port 281 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[106]
port 282 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 la_data_out[107]
port 283 nsew signal output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[108]
port 284 nsew signal output
rlabel metal2 s 154762 0 154818 800 6 la_data_out[109]
port 285 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[10]
port 286 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[110]
port 287 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[111]
port 288 nsew signal output
rlabel metal2 s 157982 0 158038 800 6 la_data_out[112]
port 289 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 la_data_out[113]
port 290 nsew signal output
rlabel metal2 s 160098 0 160154 800 6 la_data_out[114]
port 291 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 la_data_out[115]
port 292 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 la_data_out[116]
port 293 nsew signal output
rlabel metal2 s 163318 0 163374 800 6 la_data_out[117]
port 294 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 la_data_out[118]
port 295 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 la_data_out[119]
port 296 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[11]
port 297 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 la_data_out[120]
port 298 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 la_data_out[121]
port 299 nsew signal output
rlabel metal2 s 168654 0 168710 800 6 la_data_out[122]
port 300 nsew signal output
rlabel metal2 s 169758 0 169814 800 6 la_data_out[123]
port 301 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 la_data_out[124]
port 302 nsew signal output
rlabel metal2 s 171874 0 171930 800 6 la_data_out[125]
port 303 nsew signal output
rlabel metal2 s 172978 0 173034 800 6 la_data_out[126]
port 304 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 la_data_out[127]
port 305 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[12]
port 306 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[13]
port 307 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 la_data_out[14]
port 308 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[15]
port 309 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[16]
port 310 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[17]
port 311 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[18]
port 312 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[19]
port 313 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[1]
port 314 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[20]
port 315 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[21]
port 316 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[22]
port 317 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[23]
port 318 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 la_data_out[24]
port 319 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[25]
port 320 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 la_data_out[26]
port 321 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[27]
port 322 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[28]
port 323 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 la_data_out[29]
port 324 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 la_data_out[2]
port 325 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[30]
port 326 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[31]
port 327 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[32]
port 328 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[33]
port 329 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[34]
port 330 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[35]
port 331 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[36]
port 332 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[37]
port 333 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[38]
port 334 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[39]
port 335 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 la_data_out[3]
port 336 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 la_data_out[40]
port 337 nsew signal output
rlabel metal2 s 82082 0 82138 800 6 la_data_out[41]
port 338 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[42]
port 339 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[43]
port 340 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[44]
port 341 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_out[45]
port 342 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[46]
port 343 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[47]
port 344 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[48]
port 345 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[49]
port 346 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 la_data_out[4]
port 347 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[50]
port 348 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[51]
port 349 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[52]
port 350 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[53]
port 351 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[54]
port 352 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[55]
port 353 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[56]
port 354 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 la_data_out[57]
port 355 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[58]
port 356 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[59]
port 357 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[5]
port 358 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[60]
port 359 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[61]
port 360 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 la_data_out[62]
port 361 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[63]
port 362 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[64]
port 363 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[65]
port 364 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[66]
port 365 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[67]
port 366 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[68]
port 367 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[69]
port 368 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[6]
port 369 nsew signal output
rlabel metal2 s 113086 0 113142 800 6 la_data_out[70]
port 370 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[71]
port 371 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 la_data_out[72]
port 372 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 la_data_out[73]
port 373 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 la_data_out[74]
port 374 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[75]
port 375 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 la_data_out[76]
port 376 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 la_data_out[77]
port 377 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 la_data_out[78]
port 378 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 la_data_out[79]
port 379 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[7]
port 380 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[80]
port 381 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 la_data_out[81]
port 382 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 la_data_out[82]
port 383 nsew signal output
rlabel metal2 s 126978 0 127034 800 6 la_data_out[83]
port 384 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 la_data_out[84]
port 385 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 la_data_out[85]
port 386 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_out[86]
port 387 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 la_data_out[87]
port 388 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[88]
port 389 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 la_data_out[89]
port 390 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 la_data_out[8]
port 391 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[90]
port 392 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[91]
port 393 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[92]
port 394 nsew signal output
rlabel metal2 s 137650 0 137706 800 6 la_data_out[93]
port 395 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[94]
port 396 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[95]
port 397 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 la_data_out[96]
port 398 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 la_data_out[97]
port 399 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[98]
port 400 nsew signal output
rlabel metal2 s 144090 0 144146 800 6 la_data_out[99]
port 401 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[9]
port 402 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_oenb[0]
port 403 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[100]
port 404 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_oenb[101]
port 405 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 la_oenb[102]
port 406 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_oenb[103]
port 407 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_oenb[104]
port 408 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_oenb[105]
port 409 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[106]
port 410 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[107]
port 411 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oenb[108]
port 412 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oenb[109]
port 413 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_oenb[10]
port 414 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[110]
port 415 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 la_oenb[111]
port 416 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_oenb[112]
port 417 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_oenb[113]
port 418 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 la_oenb[114]
port 419 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_oenb[115]
port 420 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_oenb[116]
port 421 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_oenb[117]
port 422 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 la_oenb[118]
port 423 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_oenb[119]
port 424 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[11]
port 425 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 la_oenb[120]
port 426 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_oenb[121]
port 427 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_oenb[122]
port 428 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_oenb[123]
port 429 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_oenb[124]
port 430 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_oenb[125]
port 431 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 la_oenb[126]
port 432 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_oenb[127]
port 433 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[12]
port 434 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_oenb[13]
port 435 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[14]
port 436 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_oenb[15]
port 437 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[16]
port 438 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[17]
port 439 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[18]
port 440 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_oenb[19]
port 441 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_oenb[1]
port 442 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_oenb[20]
port 443 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[21]
port 444 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[22]
port 445 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_oenb[23]
port 446 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_oenb[24]
port 447 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[25]
port 448 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_oenb[26]
port 449 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[27]
port 450 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[28]
port 451 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oenb[29]
port 452 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[2]
port 453 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[30]
port 454 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[31]
port 455 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oenb[32]
port 456 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_oenb[33]
port 457 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[34]
port 458 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[35]
port 459 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[36]
port 460 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[37]
port 461 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[38]
port 462 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_oenb[39]
port 463 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_oenb[3]
port 464 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_oenb[40]
port 465 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_oenb[41]
port 466 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[42]
port 467 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_oenb[43]
port 468 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_oenb[44]
port 469 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[45]
port 470 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[46]
port 471 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[47]
port 472 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[48]
port 473 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_oenb[49]
port 474 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[4]
port 475 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[50]
port 476 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_oenb[51]
port 477 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[52]
port 478 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[53]
port 479 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[54]
port 480 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_oenb[55]
port 481 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_oenb[56]
port 482 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oenb[57]
port 483 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[58]
port 484 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[59]
port 485 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[5]
port 486 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_oenb[60]
port 487 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[61]
port 488 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_oenb[62]
port 489 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[63]
port 490 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[64]
port 491 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[65]
port 492 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[66]
port 493 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[67]
port 494 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[68]
port 495 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oenb[69]
port 496 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[6]
port 497 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oenb[70]
port 498 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_oenb[71]
port 499 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[72]
port 500 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_oenb[73]
port 501 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_oenb[74]
port 502 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_oenb[75]
port 503 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_oenb[76]
port 504 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_oenb[77]
port 505 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oenb[78]
port 506 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[79]
port 507 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[7]
port 508 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oenb[80]
port 509 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_oenb[81]
port 510 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_oenb[82]
port 511 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_oenb[83]
port 512 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_oenb[84]
port 513 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_oenb[85]
port 514 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_oenb[86]
port 515 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_oenb[87]
port 516 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oenb[88]
port 517 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_oenb[89]
port 518 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[8]
port 519 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[90]
port 520 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[91]
port 521 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[92]
port 522 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_oenb[93]
port 523 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[94]
port 524 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_oenb[95]
port 525 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_oenb[96]
port 526 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_oenb[97]
port 527 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_oenb[98]
port 528 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oenb[99]
port 529 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[9]
port 530 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 user_clock2
port 531 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 533 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6778518
string GDS_FILE /opt/caravel/caravel_example/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 308656
<< end >>

