magic
tech sky130A
magscale 1 2
timestamp 1647380371
<< obsli1 >>
rect 201104 202159 378848 317521
<< obsm1 >>
rect 1670 2796 583450 703044
<< metal2 >>
rect 7810 703520 7922 704960
rect 23542 703520 23654 704960
rect 39366 703520 39478 704960
rect 55098 703520 55210 704960
rect 70922 703520 71034 704960
rect 86654 703520 86766 704960
rect 102478 703520 102590 704960
rect 118210 703520 118322 704960
rect 134034 703520 134146 704960
rect 149858 703520 149970 704960
rect 165590 703520 165702 704960
rect 181414 703520 181526 704960
rect 197146 703520 197258 704960
rect 212970 703520 213082 704960
rect 228702 703520 228814 704960
rect 244526 703520 244638 704960
rect 260350 703520 260462 704960
rect 276082 703520 276194 704960
rect 291906 703520 292018 704960
rect 307638 703520 307750 704960
rect 323462 703520 323574 704960
rect 339194 703520 339306 704960
rect 355018 703520 355130 704960
rect 370842 703520 370954 704960
rect 386574 703520 386686 704960
rect 402398 703520 402510 704960
rect 418130 703520 418242 704960
rect 433954 703520 434066 704960
rect 449686 703520 449798 704960
rect 465510 703520 465622 704960
rect 481334 703520 481446 704960
rect 497066 703520 497178 704960
rect 512890 703520 513002 704960
rect 528622 703520 528734 704960
rect 544446 703520 544558 704960
rect 560178 703520 560290 704960
rect 576002 703520 576114 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17102 -960 17214 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25382 -960 25494 480
rect 26578 -960 26690 480
rect 27774 -960 27886 480
rect 28970 -960 29082 480
rect 30166 -960 30278 480
rect 31362 -960 31474 480
rect 32558 -960 32670 480
rect 33754 -960 33866 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37250 -960 37362 480
rect 38446 -960 38558 480
rect 39642 -960 39754 480
rect 40838 -960 40950 480
rect 42034 -960 42146 480
rect 43230 -960 43342 480
rect 44426 -960 44538 480
rect 45622 -960 45734 480
rect 46818 -960 46930 480
rect 48014 -960 48126 480
rect 49210 -960 49322 480
rect 50314 -960 50426 480
rect 51510 -960 51622 480
rect 52706 -960 52818 480
rect 53902 -960 54014 480
rect 55098 -960 55210 480
rect 56294 -960 56406 480
rect 57490 -960 57602 480
rect 58686 -960 58798 480
rect 59882 -960 59994 480
rect 61078 -960 61190 480
rect 62182 -960 62294 480
rect 63378 -960 63490 480
rect 64574 -960 64686 480
rect 65770 -960 65882 480
rect 66966 -960 67078 480
rect 68162 -960 68274 480
rect 69358 -960 69470 480
rect 70554 -960 70666 480
rect 71750 -960 71862 480
rect 72946 -960 73058 480
rect 74050 -960 74162 480
rect 75246 -960 75358 480
rect 76442 -960 76554 480
rect 77638 -960 77750 480
rect 78834 -960 78946 480
rect 80030 -960 80142 480
rect 81226 -960 81338 480
rect 82422 -960 82534 480
rect 83618 -960 83730 480
rect 84814 -960 84926 480
rect 85918 -960 86030 480
rect 87114 -960 87226 480
rect 88310 -960 88422 480
rect 89506 -960 89618 480
rect 90702 -960 90814 480
rect 91898 -960 92010 480
rect 93094 -960 93206 480
rect 94290 -960 94402 480
rect 95486 -960 95598 480
rect 96682 -960 96794 480
rect 97878 -960 97990 480
rect 98982 -960 99094 480
rect 100178 -960 100290 480
rect 101374 -960 101486 480
rect 102570 -960 102682 480
rect 103766 -960 103878 480
rect 104962 -960 105074 480
rect 106158 -960 106270 480
rect 107354 -960 107466 480
rect 108550 -960 108662 480
rect 109746 -960 109858 480
rect 110850 -960 110962 480
rect 112046 -960 112158 480
rect 113242 -960 113354 480
rect 114438 -960 114550 480
rect 115634 -960 115746 480
rect 116830 -960 116942 480
rect 118026 -960 118138 480
rect 119222 -960 119334 480
rect 120418 -960 120530 480
rect 121614 -960 121726 480
rect 122718 -960 122830 480
rect 123914 -960 124026 480
rect 125110 -960 125222 480
rect 126306 -960 126418 480
rect 127502 -960 127614 480
rect 128698 -960 128810 480
rect 129894 -960 130006 480
rect 131090 -960 131202 480
rect 132286 -960 132398 480
rect 133482 -960 133594 480
rect 134586 -960 134698 480
rect 135782 -960 135894 480
rect 136978 -960 137090 480
rect 138174 -960 138286 480
rect 139370 -960 139482 480
rect 140566 -960 140678 480
rect 141762 -960 141874 480
rect 142958 -960 143070 480
rect 144154 -960 144266 480
rect 145350 -960 145462 480
rect 146546 -960 146658 480
rect 147650 -960 147762 480
rect 148846 -960 148958 480
rect 150042 -960 150154 480
rect 151238 -960 151350 480
rect 152434 -960 152546 480
rect 153630 -960 153742 480
rect 154826 -960 154938 480
rect 156022 -960 156134 480
rect 157218 -960 157330 480
rect 158414 -960 158526 480
rect 159518 -960 159630 480
rect 160714 -960 160826 480
rect 161910 -960 162022 480
rect 163106 -960 163218 480
rect 164302 -960 164414 480
rect 165498 -960 165610 480
rect 166694 -960 166806 480
rect 167890 -960 168002 480
rect 169086 -960 169198 480
rect 170282 -960 170394 480
rect 171386 -960 171498 480
rect 172582 -960 172694 480
rect 173778 -960 173890 480
rect 174974 -960 175086 480
rect 176170 -960 176282 480
rect 177366 -960 177478 480
rect 178562 -960 178674 480
rect 179758 -960 179870 480
rect 180954 -960 181066 480
rect 182150 -960 182262 480
rect 183254 -960 183366 480
rect 184450 -960 184562 480
rect 185646 -960 185758 480
rect 186842 -960 186954 480
rect 188038 -960 188150 480
rect 189234 -960 189346 480
rect 190430 -960 190542 480
rect 191626 -960 191738 480
rect 192822 -960 192934 480
rect 194018 -960 194130 480
rect 195214 -960 195326 480
rect 196318 -960 196430 480
rect 197514 -960 197626 480
rect 198710 -960 198822 480
rect 199906 -960 200018 480
rect 201102 -960 201214 480
rect 202298 -960 202410 480
rect 203494 -960 203606 480
rect 204690 -960 204802 480
rect 205886 -960 205998 480
rect 207082 -960 207194 480
rect 208186 -960 208298 480
rect 209382 -960 209494 480
rect 210578 -960 210690 480
rect 211774 -960 211886 480
rect 212970 -960 213082 480
rect 214166 -960 214278 480
rect 215362 -960 215474 480
rect 216558 -960 216670 480
rect 217754 -960 217866 480
rect 218950 -960 219062 480
rect 220054 -960 220166 480
rect 221250 -960 221362 480
rect 222446 -960 222558 480
rect 223642 -960 223754 480
rect 224838 -960 224950 480
rect 226034 -960 226146 480
rect 227230 -960 227342 480
rect 228426 -960 228538 480
rect 229622 -960 229734 480
rect 230818 -960 230930 480
rect 231922 -960 232034 480
rect 233118 -960 233230 480
rect 234314 -960 234426 480
rect 235510 -960 235622 480
rect 236706 -960 236818 480
rect 237902 -960 238014 480
rect 239098 -960 239210 480
rect 240294 -960 240406 480
rect 241490 -960 241602 480
rect 242686 -960 242798 480
rect 243882 -960 243994 480
rect 244986 -960 245098 480
rect 246182 -960 246294 480
rect 247378 -960 247490 480
rect 248574 -960 248686 480
rect 249770 -960 249882 480
rect 250966 -960 251078 480
rect 252162 -960 252274 480
rect 253358 -960 253470 480
rect 254554 -960 254666 480
rect 255750 -960 255862 480
rect 256854 -960 256966 480
rect 258050 -960 258162 480
rect 259246 -960 259358 480
rect 260442 -960 260554 480
rect 261638 -960 261750 480
rect 262834 -960 262946 480
rect 264030 -960 264142 480
rect 265226 -960 265338 480
rect 266422 -960 266534 480
rect 267618 -960 267730 480
rect 268722 -960 268834 480
rect 269918 -960 270030 480
rect 271114 -960 271226 480
rect 272310 -960 272422 480
rect 273506 -960 273618 480
rect 274702 -960 274814 480
rect 275898 -960 276010 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280590 -960 280702 480
rect 281786 -960 281898 480
rect 282982 -960 283094 480
rect 284178 -960 284290 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300830 -960 300942 480
rect 302026 -960 302138 480
rect 303222 -960 303334 480
rect 304418 -960 304530 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309110 -960 309222 480
rect 310306 -960 310418 480
rect 311502 -960 311614 480
rect 312698 -960 312810 480
rect 313894 -960 314006 480
rect 315090 -960 315202 480
rect 316286 -960 316398 480
rect 317390 -960 317502 480
rect 318586 -960 318698 480
rect 319782 -960 319894 480
rect 320978 -960 321090 480
rect 322174 -960 322286 480
rect 323370 -960 323482 480
rect 324566 -960 324678 480
rect 325762 -960 325874 480
rect 326958 -960 327070 480
rect 328154 -960 328266 480
rect 329258 -960 329370 480
rect 330454 -960 330566 480
rect 331650 -960 331762 480
rect 332846 -960 332958 480
rect 334042 -960 334154 480
rect 335238 -960 335350 480
rect 336434 -960 336546 480
rect 337630 -960 337742 480
rect 338826 -960 338938 480
rect 340022 -960 340134 480
rect 341218 -960 341330 480
rect 342322 -960 342434 480
rect 343518 -960 343630 480
rect 344714 -960 344826 480
rect 345910 -960 346022 480
rect 347106 -960 347218 480
rect 348302 -960 348414 480
rect 349498 -960 349610 480
rect 350694 -960 350806 480
rect 351890 -960 352002 480
rect 353086 -960 353198 480
rect 354190 -960 354302 480
rect 355386 -960 355498 480
rect 356582 -960 356694 480
rect 357778 -960 357890 480
rect 358974 -960 359086 480
rect 360170 -960 360282 480
rect 361366 -960 361478 480
rect 362562 -960 362674 480
rect 363758 -960 363870 480
rect 364954 -960 365066 480
rect 366058 -960 366170 480
rect 367254 -960 367366 480
rect 368450 -960 368562 480
rect 369646 -960 369758 480
rect 370842 -960 370954 480
rect 372038 -960 372150 480
rect 373234 -960 373346 480
rect 374430 -960 374542 480
rect 375626 -960 375738 480
rect 376822 -960 376934 480
rect 377926 -960 378038 480
rect 379122 -960 379234 480
rect 380318 -960 380430 480
rect 381514 -960 381626 480
rect 382710 -960 382822 480
rect 383906 -960 384018 480
rect 385102 -960 385214 480
rect 386298 -960 386410 480
rect 387494 -960 387606 480
rect 388690 -960 388802 480
rect 389886 -960 389998 480
rect 390990 -960 391102 480
rect 392186 -960 392298 480
rect 393382 -960 393494 480
rect 394578 -960 394690 480
rect 395774 -960 395886 480
rect 396970 -960 397082 480
rect 398166 -960 398278 480
rect 399362 -960 399474 480
rect 400558 -960 400670 480
rect 401754 -960 401866 480
rect 402858 -960 402970 480
rect 404054 -960 404166 480
rect 405250 -960 405362 480
rect 406446 -960 406558 480
rect 407642 -960 407754 480
rect 408838 -960 408950 480
rect 410034 -960 410146 480
rect 411230 -960 411342 480
rect 412426 -960 412538 480
rect 413622 -960 413734 480
rect 414726 -960 414838 480
rect 415922 -960 416034 480
rect 417118 -960 417230 480
rect 418314 -960 418426 480
rect 419510 -960 419622 480
rect 420706 -960 420818 480
rect 421902 -960 422014 480
rect 423098 -960 423210 480
rect 424294 -960 424406 480
rect 425490 -960 425602 480
rect 426594 -960 426706 480
rect 427790 -960 427902 480
rect 428986 -960 429098 480
rect 430182 -960 430294 480
rect 431378 -960 431490 480
rect 432574 -960 432686 480
rect 433770 -960 433882 480
rect 434966 -960 435078 480
rect 436162 -960 436274 480
rect 437358 -960 437470 480
rect 438554 -960 438666 480
rect 439658 -960 439770 480
rect 440854 -960 440966 480
rect 442050 -960 442162 480
rect 443246 -960 443358 480
rect 444442 -960 444554 480
rect 445638 -960 445750 480
rect 446834 -960 446946 480
rect 448030 -960 448142 480
rect 449226 -960 449338 480
rect 450422 -960 450534 480
rect 451526 -960 451638 480
rect 452722 -960 452834 480
rect 453918 -960 454030 480
rect 455114 -960 455226 480
rect 456310 -960 456422 480
rect 457506 -960 457618 480
rect 458702 -960 458814 480
rect 459898 -960 460010 480
rect 461094 -960 461206 480
rect 462290 -960 462402 480
rect 463394 -960 463506 480
rect 464590 -960 464702 480
rect 465786 -960 465898 480
rect 466982 -960 467094 480
rect 468178 -960 468290 480
rect 469374 -960 469486 480
rect 470570 -960 470682 480
rect 471766 -960 471878 480
rect 472962 -960 473074 480
rect 474158 -960 474270 480
rect 475262 -960 475374 480
rect 476458 -960 476570 480
rect 477654 -960 477766 480
rect 478850 -960 478962 480
rect 480046 -960 480158 480
rect 481242 -960 481354 480
rect 482438 -960 482550 480
rect 483634 -960 483746 480
rect 484830 -960 484942 480
rect 486026 -960 486138 480
rect 487222 -960 487334 480
rect 488326 -960 488438 480
rect 489522 -960 489634 480
rect 490718 -960 490830 480
rect 491914 -960 492026 480
rect 493110 -960 493222 480
rect 494306 -960 494418 480
rect 495502 -960 495614 480
rect 496698 -960 496810 480
rect 497894 -960 498006 480
rect 499090 -960 499202 480
rect 500194 -960 500306 480
rect 501390 -960 501502 480
rect 502586 -960 502698 480
rect 503782 -960 503894 480
rect 504978 -960 505090 480
rect 506174 -960 506286 480
rect 507370 -960 507482 480
rect 508566 -960 508678 480
rect 509762 -960 509874 480
rect 510958 -960 511070 480
rect 512062 -960 512174 480
rect 513258 -960 513370 480
rect 514454 -960 514566 480
rect 515650 -960 515762 480
rect 516846 -960 516958 480
rect 518042 -960 518154 480
rect 519238 -960 519350 480
rect 520434 -960 520546 480
rect 521630 -960 521742 480
rect 522826 -960 522938 480
rect 523930 -960 524042 480
rect 525126 -960 525238 480
rect 526322 -960 526434 480
rect 527518 -960 527630 480
rect 528714 -960 528826 480
rect 529910 -960 530022 480
rect 531106 -960 531218 480
rect 532302 -960 532414 480
rect 533498 -960 533610 480
rect 534694 -960 534806 480
rect 535890 -960 536002 480
rect 536994 -960 537106 480
rect 538190 -960 538302 480
rect 539386 -960 539498 480
rect 540582 -960 540694 480
rect 541778 -960 541890 480
rect 542974 -960 543086 480
rect 544170 -960 544282 480
rect 545366 -960 545478 480
rect 546562 -960 546674 480
rect 547758 -960 547870 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551254 -960 551366 480
rect 552450 -960 552562 480
rect 553646 -960 553758 480
rect 554842 -960 554954 480
rect 556038 -960 556150 480
rect 557234 -960 557346 480
rect 558430 -960 558542 480
rect 559626 -960 559738 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567906 -960 568018 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 1676 703464 7754 703610
rect 7978 703464 23486 703610
rect 23710 703464 39310 703610
rect 39534 703464 55042 703610
rect 55266 703464 70866 703610
rect 71090 703464 86598 703610
rect 86822 703464 102422 703610
rect 102646 703464 118154 703610
rect 118378 703464 133978 703610
rect 134202 703464 149802 703610
rect 150026 703464 165534 703610
rect 165758 703464 181358 703610
rect 181582 703464 197090 703610
rect 197314 703464 212914 703610
rect 213138 703464 228646 703610
rect 228870 703464 244470 703610
rect 244694 703464 260294 703610
rect 260518 703464 276026 703610
rect 276250 703464 291850 703610
rect 292074 703464 307582 703610
rect 307806 703464 323406 703610
rect 323630 703464 339138 703610
rect 339362 703464 354962 703610
rect 355186 703464 370786 703610
rect 371010 703464 386518 703610
rect 386742 703464 402342 703610
rect 402566 703464 418074 703610
rect 418298 703464 433898 703610
rect 434122 703464 449630 703610
rect 449854 703464 465454 703610
rect 465678 703464 481278 703610
rect 481502 703464 497010 703610
rect 497234 703464 512834 703610
rect 513058 703464 528566 703610
rect 528790 703464 544390 703610
rect 544614 703464 560122 703610
rect 560346 703464 575946 703610
rect 576170 703464 583444 703610
rect 1676 536 583444 703464
rect 1814 326 2786 536
rect 3010 326 3982 536
rect 4206 326 5178 536
rect 5402 326 6374 536
rect 6598 326 7570 536
rect 7794 326 8766 536
rect 8990 326 9962 536
rect 10186 326 11158 536
rect 11382 326 12354 536
rect 12578 326 13458 536
rect 13682 326 14654 536
rect 14878 326 15850 536
rect 16074 326 17046 536
rect 17270 326 18242 536
rect 18466 326 19438 536
rect 19662 326 20634 536
rect 20858 326 21830 536
rect 22054 326 23026 536
rect 23250 326 24222 536
rect 24446 326 25326 536
rect 25550 326 26522 536
rect 26746 326 27718 536
rect 27942 326 28914 536
rect 29138 326 30110 536
rect 30334 326 31306 536
rect 31530 326 32502 536
rect 32726 326 33698 536
rect 33922 326 34894 536
rect 35118 326 36090 536
rect 36314 326 37194 536
rect 37418 326 38390 536
rect 38614 326 39586 536
rect 39810 326 40782 536
rect 41006 326 41978 536
rect 42202 326 43174 536
rect 43398 326 44370 536
rect 44594 326 45566 536
rect 45790 326 46762 536
rect 46986 326 47958 536
rect 48182 326 49154 536
rect 49378 326 50258 536
rect 50482 326 51454 536
rect 51678 326 52650 536
rect 52874 326 53846 536
rect 54070 326 55042 536
rect 55266 326 56238 536
rect 56462 326 57434 536
rect 57658 326 58630 536
rect 58854 326 59826 536
rect 60050 326 61022 536
rect 61246 326 62126 536
rect 62350 326 63322 536
rect 63546 326 64518 536
rect 64742 326 65714 536
rect 65938 326 66910 536
rect 67134 326 68106 536
rect 68330 326 69302 536
rect 69526 326 70498 536
rect 70722 326 71694 536
rect 71918 326 72890 536
rect 73114 326 73994 536
rect 74218 326 75190 536
rect 75414 326 76386 536
rect 76610 326 77582 536
rect 77806 326 78778 536
rect 79002 326 79974 536
rect 80198 326 81170 536
rect 81394 326 82366 536
rect 82590 326 83562 536
rect 83786 326 84758 536
rect 84982 326 85862 536
rect 86086 326 87058 536
rect 87282 326 88254 536
rect 88478 326 89450 536
rect 89674 326 90646 536
rect 90870 326 91842 536
rect 92066 326 93038 536
rect 93262 326 94234 536
rect 94458 326 95430 536
rect 95654 326 96626 536
rect 96850 326 97822 536
rect 98046 326 98926 536
rect 99150 326 100122 536
rect 100346 326 101318 536
rect 101542 326 102514 536
rect 102738 326 103710 536
rect 103934 326 104906 536
rect 105130 326 106102 536
rect 106326 326 107298 536
rect 107522 326 108494 536
rect 108718 326 109690 536
rect 109914 326 110794 536
rect 111018 326 111990 536
rect 112214 326 113186 536
rect 113410 326 114382 536
rect 114606 326 115578 536
rect 115802 326 116774 536
rect 116998 326 117970 536
rect 118194 326 119166 536
rect 119390 326 120362 536
rect 120586 326 121558 536
rect 121782 326 122662 536
rect 122886 326 123858 536
rect 124082 326 125054 536
rect 125278 326 126250 536
rect 126474 326 127446 536
rect 127670 326 128642 536
rect 128866 326 129838 536
rect 130062 326 131034 536
rect 131258 326 132230 536
rect 132454 326 133426 536
rect 133650 326 134530 536
rect 134754 326 135726 536
rect 135950 326 136922 536
rect 137146 326 138118 536
rect 138342 326 139314 536
rect 139538 326 140510 536
rect 140734 326 141706 536
rect 141930 326 142902 536
rect 143126 326 144098 536
rect 144322 326 145294 536
rect 145518 326 146490 536
rect 146714 326 147594 536
rect 147818 326 148790 536
rect 149014 326 149986 536
rect 150210 326 151182 536
rect 151406 326 152378 536
rect 152602 326 153574 536
rect 153798 326 154770 536
rect 154994 326 155966 536
rect 156190 326 157162 536
rect 157386 326 158358 536
rect 158582 326 159462 536
rect 159686 326 160658 536
rect 160882 326 161854 536
rect 162078 326 163050 536
rect 163274 326 164246 536
rect 164470 326 165442 536
rect 165666 326 166638 536
rect 166862 326 167834 536
rect 168058 326 169030 536
rect 169254 326 170226 536
rect 170450 326 171330 536
rect 171554 326 172526 536
rect 172750 326 173722 536
rect 173946 326 174918 536
rect 175142 326 176114 536
rect 176338 326 177310 536
rect 177534 326 178506 536
rect 178730 326 179702 536
rect 179926 326 180898 536
rect 181122 326 182094 536
rect 182318 326 183198 536
rect 183422 326 184394 536
rect 184618 326 185590 536
rect 185814 326 186786 536
rect 187010 326 187982 536
rect 188206 326 189178 536
rect 189402 326 190374 536
rect 190598 326 191570 536
rect 191794 326 192766 536
rect 192990 326 193962 536
rect 194186 326 195158 536
rect 195382 326 196262 536
rect 196486 326 197458 536
rect 197682 326 198654 536
rect 198878 326 199850 536
rect 200074 326 201046 536
rect 201270 326 202242 536
rect 202466 326 203438 536
rect 203662 326 204634 536
rect 204858 326 205830 536
rect 206054 326 207026 536
rect 207250 326 208130 536
rect 208354 326 209326 536
rect 209550 326 210522 536
rect 210746 326 211718 536
rect 211942 326 212914 536
rect 213138 326 214110 536
rect 214334 326 215306 536
rect 215530 326 216502 536
rect 216726 326 217698 536
rect 217922 326 218894 536
rect 219118 326 219998 536
rect 220222 326 221194 536
rect 221418 326 222390 536
rect 222614 326 223586 536
rect 223810 326 224782 536
rect 225006 326 225978 536
rect 226202 326 227174 536
rect 227398 326 228370 536
rect 228594 326 229566 536
rect 229790 326 230762 536
rect 230986 326 231866 536
rect 232090 326 233062 536
rect 233286 326 234258 536
rect 234482 326 235454 536
rect 235678 326 236650 536
rect 236874 326 237846 536
rect 238070 326 239042 536
rect 239266 326 240238 536
rect 240462 326 241434 536
rect 241658 326 242630 536
rect 242854 326 243826 536
rect 244050 326 244930 536
rect 245154 326 246126 536
rect 246350 326 247322 536
rect 247546 326 248518 536
rect 248742 326 249714 536
rect 249938 326 250910 536
rect 251134 326 252106 536
rect 252330 326 253302 536
rect 253526 326 254498 536
rect 254722 326 255694 536
rect 255918 326 256798 536
rect 257022 326 257994 536
rect 258218 326 259190 536
rect 259414 326 260386 536
rect 260610 326 261582 536
rect 261806 326 262778 536
rect 263002 326 263974 536
rect 264198 326 265170 536
rect 265394 326 266366 536
rect 266590 326 267562 536
rect 267786 326 268666 536
rect 268890 326 269862 536
rect 270086 326 271058 536
rect 271282 326 272254 536
rect 272478 326 273450 536
rect 273674 326 274646 536
rect 274870 326 275842 536
rect 276066 326 277038 536
rect 277262 326 278234 536
rect 278458 326 279430 536
rect 279654 326 280534 536
rect 280758 326 281730 536
rect 281954 326 282926 536
rect 283150 326 284122 536
rect 284346 326 285318 536
rect 285542 326 286514 536
rect 286738 326 287710 536
rect 287934 326 288906 536
rect 289130 326 290102 536
rect 290326 326 291298 536
rect 291522 326 292494 536
rect 292718 326 293598 536
rect 293822 326 294794 536
rect 295018 326 295990 536
rect 296214 326 297186 536
rect 297410 326 298382 536
rect 298606 326 299578 536
rect 299802 326 300774 536
rect 300998 326 301970 536
rect 302194 326 303166 536
rect 303390 326 304362 536
rect 304586 326 305466 536
rect 305690 326 306662 536
rect 306886 326 307858 536
rect 308082 326 309054 536
rect 309278 326 310250 536
rect 310474 326 311446 536
rect 311670 326 312642 536
rect 312866 326 313838 536
rect 314062 326 315034 536
rect 315258 326 316230 536
rect 316454 326 317334 536
rect 317558 326 318530 536
rect 318754 326 319726 536
rect 319950 326 320922 536
rect 321146 326 322118 536
rect 322342 326 323314 536
rect 323538 326 324510 536
rect 324734 326 325706 536
rect 325930 326 326902 536
rect 327126 326 328098 536
rect 328322 326 329202 536
rect 329426 326 330398 536
rect 330622 326 331594 536
rect 331818 326 332790 536
rect 333014 326 333986 536
rect 334210 326 335182 536
rect 335406 326 336378 536
rect 336602 326 337574 536
rect 337798 326 338770 536
rect 338994 326 339966 536
rect 340190 326 341162 536
rect 341386 326 342266 536
rect 342490 326 343462 536
rect 343686 326 344658 536
rect 344882 326 345854 536
rect 346078 326 347050 536
rect 347274 326 348246 536
rect 348470 326 349442 536
rect 349666 326 350638 536
rect 350862 326 351834 536
rect 352058 326 353030 536
rect 353254 326 354134 536
rect 354358 326 355330 536
rect 355554 326 356526 536
rect 356750 326 357722 536
rect 357946 326 358918 536
rect 359142 326 360114 536
rect 360338 326 361310 536
rect 361534 326 362506 536
rect 362730 326 363702 536
rect 363926 326 364898 536
rect 365122 326 366002 536
rect 366226 326 367198 536
rect 367422 326 368394 536
rect 368618 326 369590 536
rect 369814 326 370786 536
rect 371010 326 371982 536
rect 372206 326 373178 536
rect 373402 326 374374 536
rect 374598 326 375570 536
rect 375794 326 376766 536
rect 376990 326 377870 536
rect 378094 326 379066 536
rect 379290 326 380262 536
rect 380486 326 381458 536
rect 381682 326 382654 536
rect 382878 326 383850 536
rect 384074 326 385046 536
rect 385270 326 386242 536
rect 386466 326 387438 536
rect 387662 326 388634 536
rect 388858 326 389830 536
rect 390054 326 390934 536
rect 391158 326 392130 536
rect 392354 326 393326 536
rect 393550 326 394522 536
rect 394746 326 395718 536
rect 395942 326 396914 536
rect 397138 326 398110 536
rect 398334 326 399306 536
rect 399530 326 400502 536
rect 400726 326 401698 536
rect 401922 326 402802 536
rect 403026 326 403998 536
rect 404222 326 405194 536
rect 405418 326 406390 536
rect 406614 326 407586 536
rect 407810 326 408782 536
rect 409006 326 409978 536
rect 410202 326 411174 536
rect 411398 326 412370 536
rect 412594 326 413566 536
rect 413790 326 414670 536
rect 414894 326 415866 536
rect 416090 326 417062 536
rect 417286 326 418258 536
rect 418482 326 419454 536
rect 419678 326 420650 536
rect 420874 326 421846 536
rect 422070 326 423042 536
rect 423266 326 424238 536
rect 424462 326 425434 536
rect 425658 326 426538 536
rect 426762 326 427734 536
rect 427958 326 428930 536
rect 429154 326 430126 536
rect 430350 326 431322 536
rect 431546 326 432518 536
rect 432742 326 433714 536
rect 433938 326 434910 536
rect 435134 326 436106 536
rect 436330 326 437302 536
rect 437526 326 438498 536
rect 438722 326 439602 536
rect 439826 326 440798 536
rect 441022 326 441994 536
rect 442218 326 443190 536
rect 443414 326 444386 536
rect 444610 326 445582 536
rect 445806 326 446778 536
rect 447002 326 447974 536
rect 448198 326 449170 536
rect 449394 326 450366 536
rect 450590 326 451470 536
rect 451694 326 452666 536
rect 452890 326 453862 536
rect 454086 326 455058 536
rect 455282 326 456254 536
rect 456478 326 457450 536
rect 457674 326 458646 536
rect 458870 326 459842 536
rect 460066 326 461038 536
rect 461262 326 462234 536
rect 462458 326 463338 536
rect 463562 326 464534 536
rect 464758 326 465730 536
rect 465954 326 466926 536
rect 467150 326 468122 536
rect 468346 326 469318 536
rect 469542 326 470514 536
rect 470738 326 471710 536
rect 471934 326 472906 536
rect 473130 326 474102 536
rect 474326 326 475206 536
rect 475430 326 476402 536
rect 476626 326 477598 536
rect 477822 326 478794 536
rect 479018 326 479990 536
rect 480214 326 481186 536
rect 481410 326 482382 536
rect 482606 326 483578 536
rect 483802 326 484774 536
rect 484998 326 485970 536
rect 486194 326 487166 536
rect 487390 326 488270 536
rect 488494 326 489466 536
rect 489690 326 490662 536
rect 490886 326 491858 536
rect 492082 326 493054 536
rect 493278 326 494250 536
rect 494474 326 495446 536
rect 495670 326 496642 536
rect 496866 326 497838 536
rect 498062 326 499034 536
rect 499258 326 500138 536
rect 500362 326 501334 536
rect 501558 326 502530 536
rect 502754 326 503726 536
rect 503950 326 504922 536
rect 505146 326 506118 536
rect 506342 326 507314 536
rect 507538 326 508510 536
rect 508734 326 509706 536
rect 509930 326 510902 536
rect 511126 326 512006 536
rect 512230 326 513202 536
rect 513426 326 514398 536
rect 514622 326 515594 536
rect 515818 326 516790 536
rect 517014 326 517986 536
rect 518210 326 519182 536
rect 519406 326 520378 536
rect 520602 326 521574 536
rect 521798 326 522770 536
rect 522994 326 523874 536
rect 524098 326 525070 536
rect 525294 326 526266 536
rect 526490 326 527462 536
rect 527686 326 528658 536
rect 528882 326 529854 536
rect 530078 326 531050 536
rect 531274 326 532246 536
rect 532470 326 533442 536
rect 533666 326 534638 536
rect 534862 326 535834 536
rect 536058 326 536938 536
rect 537162 326 538134 536
rect 538358 326 539330 536
rect 539554 326 540526 536
rect 540750 326 541722 536
rect 541946 326 542918 536
rect 543142 326 544114 536
rect 544338 326 545310 536
rect 545534 326 546506 536
rect 546730 326 547702 536
rect 547926 326 548806 536
rect 549030 326 550002 536
rect 550226 326 551198 536
rect 551422 326 552394 536
rect 552618 326 553590 536
rect 553814 326 554786 536
rect 555010 326 555982 536
rect 556206 326 557178 536
rect 557402 326 558374 536
rect 558598 326 559570 536
rect 559794 326 560674 536
rect 560898 326 561870 536
rect 562094 326 563066 536
rect 563290 326 564262 536
rect 564486 326 565458 536
rect 565682 326 566654 536
rect 566878 326 567850 536
rect 568074 326 569046 536
rect 569270 326 570242 536
rect 570466 326 571438 536
rect 571662 326 572542 536
rect 572766 326 573738 536
rect 573962 326 574934 536
rect 575158 326 576130 536
rect 576354 326 577326 536
rect 577550 326 578522 536
rect 578746 326 579718 536
rect 579942 326 580914 536
rect 581138 326 582110 536
rect 582334 326 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697220 584960 697460
rect -960 684164 480 684404
rect 583520 684164 584960 684404
rect -960 671108 480 671348
rect 583520 671108 584960 671348
rect -960 658052 480 658292
rect 583520 658052 584960 658292
rect -960 644996 480 645236
rect 583520 644996 584960 645236
rect -960 631940 480 632180
rect 583520 631940 584960 632180
rect -960 619020 480 619260
rect 583520 619020 584960 619260
rect -960 605964 480 606204
rect 583520 605964 584960 606204
rect -960 592908 480 593148
rect 583520 592908 584960 593148
rect -960 579852 480 580092
rect 583520 579852 584960 580092
rect -960 566796 480 567036
rect 583520 566796 584960 567036
rect -960 553740 480 553980
rect 583520 553740 584960 553980
rect -960 540684 480 540924
rect 583520 540684 584960 540924
rect -960 527764 480 528004
rect 583520 527764 584960 528004
rect -960 514708 480 514948
rect 583520 514708 584960 514948
rect -960 501652 480 501892
rect 583520 501652 584960 501892
rect -960 488596 480 488836
rect 583520 488596 584960 488836
rect -960 475540 480 475780
rect 583520 475540 584960 475780
rect -960 462484 480 462724
rect 583520 462484 584960 462724
rect -960 449428 480 449668
rect 583520 449428 584960 449668
rect -960 436508 480 436748
rect 583520 436508 584960 436748
rect -960 423452 480 423692
rect 583520 423452 584960 423692
rect -960 410396 480 410636
rect 583520 410396 584960 410636
rect -960 397340 480 397580
rect 583520 397340 584960 397580
rect -960 384284 480 384524
rect 583520 384284 584960 384524
rect -960 371228 480 371468
rect 583520 371228 584960 371468
rect -960 358308 480 358548
rect 583520 358308 584960 358548
rect -960 345252 480 345492
rect 583520 345252 584960 345492
rect -960 332196 480 332436
rect 583520 332196 584960 332436
rect -960 319140 480 319380
rect 583520 319140 584960 319380
rect -960 306084 480 306324
rect 583520 306084 584960 306324
rect -960 293028 480 293268
rect 583520 293028 584960 293268
rect -960 279972 480 280212
rect 583520 279972 584960 280212
rect -960 267052 480 267292
rect 583520 267052 584960 267292
rect -960 253996 480 254236
rect 583520 253996 584960 254236
rect -960 240940 480 241180
rect 583520 240940 584960 241180
rect -960 227884 480 228124
rect 583520 227884 584960 228124
rect -960 214828 480 215068
rect 583520 214828 584960 215068
rect -960 201772 480 202012
rect 583520 201772 584960 202012
rect -960 188716 480 188956
rect 583520 188716 584960 188956
rect -960 175796 480 176036
rect 583520 175796 584960 176036
rect -960 162740 480 162980
rect 583520 162740 584960 162980
rect -960 149684 480 149924
rect 583520 149684 584960 149924
rect -960 136628 480 136868
rect 583520 136628 584960 136868
rect -960 123572 480 123812
rect 583520 123572 584960 123812
rect -960 110516 480 110756
rect 583520 110516 584960 110756
rect -960 97460 480 97700
rect 583520 97460 584960 97700
rect -960 84540 480 84780
rect 583520 84540 584960 84780
rect -960 71484 480 71724
rect 583520 71484 584960 71724
rect -960 58428 480 58668
rect 583520 58428 584960 58668
rect -960 45372 480 45612
rect 583520 45372 584960 45612
rect -960 32316 480 32556
rect 583520 32316 584960 32556
rect -960 19260 480 19500
rect 583520 19260 584960 19500
rect -960 6340 480 6580
rect 583520 6340 584960 6580
<< obsm3 >>
rect 560 697140 583440 697373
rect 246 684484 583586 697140
rect 560 684084 583440 684484
rect 246 671428 583586 684084
rect 560 671028 583440 671428
rect 246 658372 583586 671028
rect 560 657972 583440 658372
rect 246 645316 583586 657972
rect 560 644916 583440 645316
rect 246 632260 583586 644916
rect 560 631860 583440 632260
rect 246 619340 583586 631860
rect 560 618940 583440 619340
rect 246 606284 583586 618940
rect 560 605884 583440 606284
rect 246 593228 583586 605884
rect 560 592828 583440 593228
rect 246 580172 583586 592828
rect 560 579772 583440 580172
rect 246 567116 583586 579772
rect 560 566716 583440 567116
rect 246 554060 583586 566716
rect 560 553660 583440 554060
rect 246 541004 583586 553660
rect 560 540604 583440 541004
rect 246 528084 583586 540604
rect 560 527684 583440 528084
rect 246 515028 583586 527684
rect 560 514628 583440 515028
rect 246 501972 583586 514628
rect 560 501572 583440 501972
rect 246 488916 583586 501572
rect 560 488516 583440 488916
rect 246 475860 583586 488516
rect 560 475460 583440 475860
rect 246 462804 583586 475460
rect 560 462404 583440 462804
rect 246 449748 583586 462404
rect 560 449348 583440 449748
rect 246 436828 583586 449348
rect 560 436428 583440 436828
rect 246 423772 583586 436428
rect 560 423372 583440 423772
rect 246 410716 583586 423372
rect 560 410316 583440 410716
rect 246 397660 583586 410316
rect 560 397260 583440 397660
rect 246 384604 583586 397260
rect 560 384204 583440 384604
rect 246 371548 583586 384204
rect 560 371148 583440 371548
rect 246 358628 583586 371148
rect 560 358228 583440 358628
rect 246 345572 583586 358228
rect 560 345172 583440 345572
rect 246 332516 583586 345172
rect 560 332116 583440 332516
rect 246 319460 583586 332116
rect 560 319060 583440 319460
rect 246 306404 583586 319060
rect 560 306004 583440 306404
rect 246 293348 583586 306004
rect 560 292948 583440 293348
rect 246 280292 583586 292948
rect 560 279892 583440 280292
rect 246 267372 583586 279892
rect 560 266972 583440 267372
rect 246 254316 583586 266972
rect 560 253916 583440 254316
rect 246 241260 583586 253916
rect 560 240860 583440 241260
rect 246 228204 583586 240860
rect 560 227804 583440 228204
rect 246 215148 583586 227804
rect 560 214748 583440 215148
rect 246 202092 583586 214748
rect 560 201692 583440 202092
rect 246 189036 583586 201692
rect 560 188636 583440 189036
rect 246 176116 583586 188636
rect 560 175716 583440 176116
rect 246 163060 583586 175716
rect 560 162660 583440 163060
rect 246 150004 583586 162660
rect 560 149604 583440 150004
rect 246 136948 583586 149604
rect 560 136548 583440 136948
rect 246 123892 583586 136548
rect 560 123492 583440 123892
rect 246 110836 583586 123492
rect 560 110436 583440 110836
rect 246 97780 583586 110436
rect 560 97380 583440 97780
rect 246 84860 583586 97380
rect 560 84460 583440 84860
rect 246 71804 583586 84460
rect 560 71404 583440 71804
rect 246 58748 583586 71404
rect 560 58348 583440 58748
rect 246 45692 583586 58348
rect 560 45292 583440 45692
rect 246 32636 583586 45292
rect 560 32236 583440 32636
rect 246 19580 583586 32236
rect 560 19180 583440 19580
rect 246 6660 583586 19180
rect 560 6260 583440 6660
rect 246 3299 583586 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 9234 -5734 9854 709670
rect 12954 -7654 13574 711590
rect 19794 -1894 20414 705830
rect 23514 -3814 24134 707750
rect 27234 -5734 27854 709670
rect 30954 -7654 31574 711590
rect 37794 -1894 38414 705830
rect 41514 -3814 42134 707750
rect 45234 -5734 45854 709670
rect 48954 -7654 49574 711590
rect 55794 -1894 56414 705830
rect 59514 -3814 60134 707750
rect 63234 -5734 63854 709670
rect 66954 -7654 67574 711590
rect 73794 -1894 74414 705830
rect 77514 -3814 78134 707750
rect 81234 -5734 81854 709670
rect 84954 -7654 85574 711590
rect 91794 -1894 92414 705830
rect 95514 -3814 96134 707750
rect 99234 -5734 99854 709670
rect 102954 -7654 103574 711590
rect 109794 -1894 110414 705830
rect 113514 -3814 114134 707750
rect 117234 -5734 117854 709670
rect 120954 -7654 121574 711590
rect 127794 -1894 128414 705830
rect 131514 -3814 132134 707750
rect 135234 -5734 135854 709670
rect 138954 -7654 139574 711590
rect 145794 -1894 146414 705830
rect 149514 -3814 150134 707750
rect 153234 -5734 153854 709670
rect 156954 -7654 157574 711590
rect 163794 -1894 164414 705830
rect 167514 -3814 168134 707750
rect 171234 -5734 171854 709670
rect 174954 -7654 175574 711590
rect 181794 -1894 182414 705830
rect 185514 -3814 186134 707750
rect 189234 -5734 189854 709670
rect 192954 -7654 193574 711590
rect 199794 322000 200414 705830
rect 203514 322000 204134 707750
rect 207234 322000 207854 709670
rect 210954 322000 211574 711590
rect 217794 322000 218414 705830
rect 221514 322000 222134 707750
rect 225234 322000 225854 709670
rect 228954 322000 229574 711590
rect 235794 322000 236414 705830
rect 239514 322000 240134 707750
rect 243234 322000 243854 709670
rect 246954 322000 247574 711590
rect 253794 322000 254414 705830
rect 257514 322000 258134 707750
rect 261234 322000 261854 709670
rect 264954 322000 265574 711590
rect 271794 322000 272414 705830
rect 275514 322000 276134 707750
rect 279234 322000 279854 709670
rect 282954 322000 283574 711590
rect 289794 322000 290414 705830
rect 293514 322000 294134 707750
rect 297234 322000 297854 709670
rect 300954 322000 301574 711590
rect 307794 322000 308414 705830
rect 311514 322000 312134 707750
rect 315234 322000 315854 709670
rect 318954 322000 319574 711590
rect 325794 322000 326414 705830
rect 329514 322000 330134 707750
rect 333234 322000 333854 709670
rect 336954 322000 337574 711590
rect 343794 322000 344414 705830
rect 347514 322000 348134 707750
rect 351234 322000 351854 709670
rect 354954 322000 355574 711590
rect 361794 322000 362414 705830
rect 365514 322000 366134 707750
rect 369234 322000 369854 709670
rect 372954 322000 373574 711590
rect 379794 322000 380414 705830
rect 199794 -1894 200414 198000
rect 203514 -3814 204134 198000
rect 207234 -5734 207854 198000
rect 210954 -7654 211574 198000
rect 217794 -1894 218414 198000
rect 221514 -3814 222134 198000
rect 225234 -5734 225854 198000
rect 228954 -7654 229574 198000
rect 235794 -1894 236414 198000
rect 239514 -3814 240134 198000
rect 243234 -5734 243854 198000
rect 246954 -7654 247574 198000
rect 253794 -1894 254414 198000
rect 257514 -3814 258134 198000
rect 261234 -5734 261854 198000
rect 264954 -7654 265574 198000
rect 271794 -1894 272414 198000
rect 275514 -3814 276134 198000
rect 279234 -5734 279854 198000
rect 282954 -7654 283574 198000
rect 289794 -1894 290414 198000
rect 293514 -3814 294134 198000
rect 297234 -5734 297854 198000
rect 300954 -7654 301574 198000
rect 307794 -1894 308414 198000
rect 311514 -3814 312134 198000
rect 315234 -5734 315854 198000
rect 318954 -7654 319574 198000
rect 325794 -1894 326414 198000
rect 329514 -3814 330134 198000
rect 333234 -5734 333854 198000
rect 336954 -7654 337574 198000
rect 343794 -1894 344414 198000
rect 347514 -3814 348134 198000
rect 351234 -5734 351854 198000
rect 354954 -7654 355574 198000
rect 361794 -1894 362414 198000
rect 365514 -3814 366134 198000
rect 369234 -5734 369854 198000
rect 372954 -7654 373574 198000
rect 379794 -1894 380414 198000
rect 383514 -3814 384134 707750
rect 387234 -5734 387854 709670
rect 390954 -7654 391574 711590
rect 397794 -1894 398414 705830
rect 401514 -3814 402134 707750
rect 405234 -5734 405854 709670
rect 408954 -7654 409574 711590
rect 415794 -1894 416414 705830
rect 419514 -3814 420134 707750
rect 423234 -5734 423854 709670
rect 426954 -7654 427574 711590
rect 433794 -1894 434414 705830
rect 437514 -3814 438134 707750
rect 441234 -5734 441854 709670
rect 444954 -7654 445574 711590
rect 451794 -1894 452414 705830
rect 455514 -3814 456134 707750
rect 459234 -5734 459854 709670
rect 462954 -7654 463574 711590
rect 469794 -1894 470414 705830
rect 473514 -3814 474134 707750
rect 477234 -5734 477854 709670
rect 480954 -7654 481574 711590
rect 487794 -1894 488414 705830
rect 491514 -3814 492134 707750
rect 495234 -5734 495854 709670
rect 498954 -7654 499574 711590
rect 505794 -1894 506414 705830
rect 509514 -3814 510134 707750
rect 513234 -5734 513854 709670
rect 516954 -7654 517574 711590
rect 523794 -1894 524414 705830
rect 527514 -3814 528134 707750
rect 531234 -5734 531854 709670
rect 534954 -7654 535574 711590
rect 541794 -1894 542414 705830
rect 545514 -3814 546134 707750
rect 549234 -5734 549854 709670
rect 552954 -7654 553574 711590
rect 559794 -1894 560414 705830
rect 563514 -3814 564134 707750
rect 567234 -5734 567854 709670
rect 570954 -7654 571574 711590
rect 577794 -1894 578414 705830
rect 581514 -3814 582134 707750
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 3371 6427 5434 322149
rect 6214 6427 9154 322149
rect 9934 6427 12874 322149
rect 13654 6427 19714 322149
rect 20494 6427 23434 322149
rect 24214 6427 27154 322149
rect 27934 6427 30874 322149
rect 31654 6427 37714 322149
rect 38494 6427 41434 322149
rect 42214 6427 45154 322149
rect 45934 6427 48874 322149
rect 49654 6427 55714 322149
rect 56494 6427 59434 322149
rect 60214 6427 63154 322149
rect 63934 6427 66874 322149
rect 67654 6427 73714 322149
rect 74494 6427 77434 322149
rect 78214 6427 81154 322149
rect 81934 6427 84874 322149
rect 85654 6427 91714 322149
rect 92494 6427 95434 322149
rect 96214 6427 99154 322149
rect 99934 6427 102874 322149
rect 103654 6427 109714 322149
rect 110494 6427 113434 322149
rect 114214 6427 117154 322149
rect 117934 6427 120874 322149
rect 121654 6427 127714 322149
rect 128494 6427 131434 322149
rect 132214 6427 135154 322149
rect 135934 6427 138874 322149
rect 139654 6427 145714 322149
rect 146494 6427 149434 322149
rect 150214 6427 153154 322149
rect 153934 6427 156874 322149
rect 157654 6427 163714 322149
rect 164494 6427 167434 322149
rect 168214 6427 171154 322149
rect 171934 6427 174874 322149
rect 175654 6427 181714 322149
rect 182494 6427 185434 322149
rect 186214 6427 189154 322149
rect 189934 6427 192874 322149
rect 193654 321920 199714 322149
rect 200494 321920 203434 322149
rect 204214 321920 207154 322149
rect 207934 321920 210874 322149
rect 211654 321920 217714 322149
rect 218494 321920 221434 322149
rect 222214 321920 225154 322149
rect 225934 321920 228874 322149
rect 229654 321920 235714 322149
rect 236494 321920 239434 322149
rect 240214 321920 243154 322149
rect 243934 321920 246874 322149
rect 247654 321920 253714 322149
rect 254494 321920 257434 322149
rect 258214 321920 261154 322149
rect 261934 321920 264874 322149
rect 265654 321920 271714 322149
rect 272494 321920 275434 322149
rect 276214 321920 279154 322149
rect 279934 321920 282874 322149
rect 283654 321920 289714 322149
rect 290494 321920 293434 322149
rect 294214 321920 297154 322149
rect 297934 321920 300874 322149
rect 301654 321920 307714 322149
rect 308494 321920 311434 322149
rect 312214 321920 315154 322149
rect 315934 321920 318874 322149
rect 319654 321920 325714 322149
rect 326494 321920 329434 322149
rect 330214 321920 333154 322149
rect 333934 321920 336874 322149
rect 337654 321920 343714 322149
rect 344494 321920 347434 322149
rect 348214 321920 351154 322149
rect 351934 321920 354874 322149
rect 355654 321920 361714 322149
rect 362494 321920 365434 322149
rect 366214 321920 369154 322149
rect 369934 321920 372874 322149
rect 373654 321920 379714 322149
rect 380494 321920 383434 322149
rect 193654 198080 383434 321920
rect 193654 6427 199714 198080
rect 200494 6427 203434 198080
rect 204214 6427 207154 198080
rect 207934 6427 210874 198080
rect 211654 6427 217714 198080
rect 218494 6427 221434 198080
rect 222214 6427 225154 198080
rect 225934 6427 228874 198080
rect 229654 6427 235714 198080
rect 236494 6427 239434 198080
rect 240214 6427 243154 198080
rect 243934 6427 246874 198080
rect 247654 6427 253714 198080
rect 254494 6427 257434 198080
rect 258214 6427 261154 198080
rect 261934 6427 264874 198080
rect 265654 6427 271714 198080
rect 272494 6427 275434 198080
rect 276214 6427 279154 198080
rect 279934 6427 282874 198080
rect 283654 6427 289714 198080
rect 290494 6427 293434 198080
rect 294214 6427 297154 198080
rect 297934 6427 300874 198080
rect 301654 6427 307714 198080
rect 308494 6427 311434 198080
rect 312214 6427 315154 198080
rect 315934 6427 318874 198080
rect 319654 6427 325714 198080
rect 326494 6427 329434 198080
rect 330214 6427 333154 198080
rect 333934 6427 336874 198080
rect 337654 6427 343714 198080
rect 344494 6427 347434 198080
rect 348214 6427 351154 198080
rect 351934 6427 354874 198080
rect 355654 6427 361714 198080
rect 362494 6427 365434 198080
rect 366214 6427 369154 198080
rect 369934 6427 372874 198080
rect 373654 6427 379714 198080
rect 380494 6427 383434 198080
rect 384214 6427 387154 322149
rect 387934 6427 390874 322149
rect 391654 6427 397714 322149
rect 398494 6427 401434 322149
rect 402214 6427 405154 322149
rect 405934 6427 408874 322149
rect 409654 6427 415714 322149
rect 416494 6427 419434 322149
rect 420214 6427 423154 322149
rect 423934 6427 426874 322149
rect 427654 6427 433714 322149
rect 434494 6427 437434 322149
rect 438214 6427 441154 322149
rect 441934 6427 444874 322149
rect 445654 6427 451714 322149
rect 452494 6427 455434 322149
rect 456214 6427 459154 322149
rect 459934 6427 462874 322149
rect 463654 6427 469714 322149
rect 470494 6427 473434 322149
rect 474214 6427 477154 322149
rect 477934 6427 480874 322149
rect 481654 6427 487714 322149
rect 488494 6427 491434 322149
rect 492214 6427 495154 322149
rect 495934 6427 498874 322149
rect 499654 6427 505714 322149
rect 506494 6427 509434 322149
rect 510214 6427 513154 322149
rect 513934 6427 516874 322149
rect 517654 6427 523714 322149
rect 524494 6427 527434 322149
rect 528214 6427 531154 322149
rect 531934 6427 534874 322149
rect 535654 6427 541714 322149
rect 542494 6427 545434 322149
rect 546214 6427 549154 322149
rect 549934 6427 552874 322149
rect 553654 6427 559714 322149
rect 560494 6427 563434 322149
rect 564214 6427 567154 322149
rect 567934 6427 570874 322149
rect 571654 6427 577714 322149
rect 578494 6427 580461 322149
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -6806 694306 590730 694926
rect -4886 690586 588810 691206
rect -2966 686866 586890 687486
rect -8726 680026 592650 680646
rect -6806 676306 590730 676926
rect -4886 672586 588810 673206
rect -2966 668866 586890 669486
rect -8726 662026 592650 662646
rect -6806 658306 590730 658926
rect -4886 654586 588810 655206
rect -2966 650866 586890 651486
rect -8726 644026 592650 644646
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -2966 632866 586890 633486
rect -8726 626026 592650 626646
rect -6806 622306 590730 622926
rect -4886 618586 588810 619206
rect -2966 614866 586890 615486
rect -8726 608026 592650 608646
rect -6806 604306 590730 604926
rect -4886 600586 588810 601206
rect -2966 596866 586890 597486
rect -8726 590026 592650 590646
rect -6806 586306 590730 586926
rect -4886 582586 588810 583206
rect -2966 578866 586890 579486
rect -8726 572026 592650 572646
rect -6806 568306 590730 568926
rect -4886 564586 588810 565206
rect -2966 560866 586890 561486
rect -8726 554026 592650 554646
rect -6806 550306 590730 550926
rect -4886 546586 588810 547206
rect -2966 542866 586890 543486
rect -8726 536026 592650 536646
rect -6806 532306 590730 532926
rect -4886 528586 588810 529206
rect -2966 524866 586890 525486
rect -8726 518026 592650 518646
rect -6806 514306 590730 514926
rect -4886 510586 588810 511206
rect -2966 506866 586890 507486
rect -8726 500026 592650 500646
rect -6806 496306 590730 496926
rect -4886 492586 588810 493206
rect -2966 488866 586890 489486
rect -8726 482026 592650 482646
rect -6806 478306 590730 478926
rect -4886 474586 588810 475206
rect -2966 470866 586890 471486
rect -8726 464026 592650 464646
rect -6806 460306 590730 460926
rect -4886 456586 588810 457206
rect -2966 452866 586890 453486
rect -8726 446026 592650 446646
rect -6806 442306 590730 442926
rect -4886 438586 588810 439206
rect -2966 434866 586890 435486
rect -8726 428026 592650 428646
rect -6806 424306 590730 424926
rect -4886 420586 588810 421206
rect -2966 416866 586890 417486
rect -8726 410026 592650 410646
rect -6806 406306 590730 406926
rect -4886 402586 588810 403206
rect -2966 398866 586890 399486
rect -8726 392026 592650 392646
rect -6806 388306 590730 388926
rect -4886 384586 588810 385206
rect -2966 380866 586890 381486
rect -8726 374026 592650 374646
rect -6806 370306 590730 370926
rect -4886 366586 588810 367206
rect -2966 362866 586890 363486
rect -8726 356026 592650 356646
rect -6806 352306 590730 352926
rect -4886 348586 588810 349206
rect -2966 344866 586890 345486
rect -8726 338026 592650 338646
rect -6806 334306 590730 334926
rect -4886 330586 588810 331206
rect -2966 326866 586890 327486
rect -8726 320026 592650 320646
rect -6806 316306 590730 316926
rect -4886 312586 588810 313206
rect -2966 308866 586890 309486
rect -8726 302026 592650 302646
rect -6806 298306 590730 298926
rect -4886 294586 588810 295206
rect -2966 290866 586890 291486
rect -8726 284026 592650 284646
rect -6806 280306 590730 280926
rect -4886 276586 588810 277206
rect -2966 272866 586890 273486
rect -8726 266026 592650 266646
rect -6806 262306 590730 262926
rect -4886 258586 588810 259206
rect -2966 254866 586890 255486
rect -8726 248026 592650 248646
rect -6806 244306 590730 244926
rect -4886 240586 588810 241206
rect -2966 236866 586890 237486
rect -8726 230026 592650 230646
rect -6806 226306 590730 226926
rect -4886 222586 588810 223206
rect -2966 218866 586890 219486
rect -8726 212026 592650 212646
rect -6806 208306 590730 208926
rect -4886 204586 588810 205206
rect -2966 200866 586890 201486
rect -8726 194026 592650 194646
rect -6806 190306 590730 190926
rect -4886 186586 588810 187206
rect -2966 182866 586890 183486
rect -8726 176026 592650 176646
rect -6806 172306 590730 172926
rect -4886 168586 588810 169206
rect -2966 164866 586890 165486
rect -8726 158026 592650 158646
rect -6806 154306 590730 154926
rect -4886 150586 588810 151206
rect -2966 146866 586890 147486
rect -8726 140026 592650 140646
rect -6806 136306 590730 136926
rect -4886 132586 588810 133206
rect -2966 128866 586890 129486
rect -8726 122026 592650 122646
rect -6806 118306 590730 118926
rect -4886 114586 588810 115206
rect -2966 110866 586890 111486
rect -8726 104026 592650 104646
rect -6806 100306 590730 100926
rect -4886 96586 588810 97206
rect -2966 92866 586890 93486
rect -8726 86026 592650 86646
rect -6806 82306 590730 82926
rect -4886 78586 588810 79206
rect -2966 74866 586890 75486
rect -8726 68026 592650 68646
rect -6806 64306 590730 64926
rect -4886 60586 588810 61206
rect -2966 56866 586890 57486
rect -8726 50026 592650 50646
rect -6806 46306 590730 46926
rect -4886 42586 588810 43206
rect -2966 38866 586890 39486
rect -8726 32026 592650 32646
rect -6806 28306 590730 28926
rect -4886 24586 588810 25206
rect -2966 20866 586890 21486
rect -8726 14026 592650 14646
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 279972 584960 280212 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 449686 703520 449798 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 386574 703520 386686 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 323462 703520 323574 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 260350 703520 260462 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 197146 703520 197258 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 134034 703520 134146 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 70922 703520 71034 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 332196 584960 332436 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 384284 584960 384524 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 436508 584960 436748 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 488596 584960 488836 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 540684 584960 540924 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 592908 584960 593148 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 644996 584960 645236 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 576002 703520 576114 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 512890 703520 513002 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6340 584960 6580 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 449428 584960 449668 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 501652 584960 501892 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 553740 584960 553980 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 605964 584960 606204 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 658052 584960 658292 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 560178 703520 560290 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 497066 703520 497178 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 433954 703520 434066 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 370842 703520 370954 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 307638 703520 307750 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 45372 584960 45612 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 244526 703520 244638 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 181414 703520 181526 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 118210 703520 118322 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 55098 703520 55210 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 84540 584960 84780 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 123572 584960 123812 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 162740 584960 162980 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 201772 584960 202012 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 240940 584960 241180 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 293028 584960 293268 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 345252 584960 345492 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 397340 584960 397580 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32316 584960 32556 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 475540 584960 475780 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 527764 584960 528004 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 579852 584960 580092 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 631940 584960 632180 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 684164 584960 684404 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 528622 703520 528734 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 465510 703520 465622 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 402398 703520 402510 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 339194 703520 339306 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 276082 703520 276194 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 71484 584960 71724 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 212970 703520 213082 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 149858 703520 149970 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 86654 703520 86766 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 23542 703520 23654 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 110516 584960 110756 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 149684 584960 149924 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 188716 584960 188956 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 227884 584960 228124 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 267052 584960 267292 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 319140 584960 319380 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 371228 584960 371468 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 423452 584960 423692 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19260 584960 19500 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 462484 584960 462724 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 514708 584960 514948 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 566796 584960 567036 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 619020 584960 619260 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 671108 584960 671348 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 544446 703520 544558 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 481334 703520 481446 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 418130 703520 418242 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 355018 703520 355130 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 291906 703520 292018 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 58428 584960 58668 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 228702 703520 228814 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 165590 703520 165702 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 102478 703520 102590 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 39366 703520 39478 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 97460 584960 97700 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 136628 584960 136868 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 175796 584960 176036 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 214828 584960 215068 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 253996 584960 254236 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 306084 584960 306324 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 358308 584960 358548 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 410396 584960 410636 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 irq[0]
port 144 nsew signal output
rlabel metal2 s 7810 703520 7922 704960 6 irq[1]
port 145 nsew signal output
rlabel metal3 s 583520 697220 584960 697460 6 irq[2]
port 146 nsew signal output
rlabel metal2 s 126306 -960 126418 480 8 la_data_in[0]
port 147 nsew signal input
rlabel metal2 s 482438 -960 482550 480 8 la_data_in[100]
port 148 nsew signal input
rlabel metal2 s 486026 -960 486138 480 8 la_data_in[101]
port 149 nsew signal input
rlabel metal2 s 489522 -960 489634 480 8 la_data_in[102]
port 150 nsew signal input
rlabel metal2 s 493110 -960 493222 480 8 la_data_in[103]
port 151 nsew signal input
rlabel metal2 s 496698 -960 496810 480 8 la_data_in[104]
port 152 nsew signal input
rlabel metal2 s 500194 -960 500306 480 8 la_data_in[105]
port 153 nsew signal input
rlabel metal2 s 503782 -960 503894 480 8 la_data_in[106]
port 154 nsew signal input
rlabel metal2 s 507370 -960 507482 480 8 la_data_in[107]
port 155 nsew signal input
rlabel metal2 s 510958 -960 511070 480 8 la_data_in[108]
port 156 nsew signal input
rlabel metal2 s 514454 -960 514566 480 8 la_data_in[109]
port 157 nsew signal input
rlabel metal2 s 161910 -960 162022 480 8 la_data_in[10]
port 158 nsew signal input
rlabel metal2 s 518042 -960 518154 480 8 la_data_in[110]
port 159 nsew signal input
rlabel metal2 s 521630 -960 521742 480 8 la_data_in[111]
port 160 nsew signal input
rlabel metal2 s 525126 -960 525238 480 8 la_data_in[112]
port 161 nsew signal input
rlabel metal2 s 528714 -960 528826 480 8 la_data_in[113]
port 162 nsew signal input
rlabel metal2 s 532302 -960 532414 480 8 la_data_in[114]
port 163 nsew signal input
rlabel metal2 s 535890 -960 536002 480 8 la_data_in[115]
port 164 nsew signal input
rlabel metal2 s 539386 -960 539498 480 8 la_data_in[116]
port 165 nsew signal input
rlabel metal2 s 542974 -960 543086 480 8 la_data_in[117]
port 166 nsew signal input
rlabel metal2 s 546562 -960 546674 480 8 la_data_in[118]
port 167 nsew signal input
rlabel metal2 s 550058 -960 550170 480 8 la_data_in[119]
port 168 nsew signal input
rlabel metal2 s 165498 -960 165610 480 8 la_data_in[11]
port 169 nsew signal input
rlabel metal2 s 553646 -960 553758 480 8 la_data_in[120]
port 170 nsew signal input
rlabel metal2 s 557234 -960 557346 480 8 la_data_in[121]
port 171 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 la_data_in[122]
port 172 nsew signal input
rlabel metal2 s 564318 -960 564430 480 8 la_data_in[123]
port 173 nsew signal input
rlabel metal2 s 567906 -960 568018 480 8 la_data_in[124]
port 174 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_data_in[125]
port 175 nsew signal input
rlabel metal2 s 574990 -960 575102 480 8 la_data_in[126]
port 176 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_data_in[127]
port 177 nsew signal input
rlabel metal2 s 169086 -960 169198 480 8 la_data_in[12]
port 178 nsew signal input
rlabel metal2 s 172582 -960 172694 480 8 la_data_in[13]
port 179 nsew signal input
rlabel metal2 s 176170 -960 176282 480 8 la_data_in[14]
port 180 nsew signal input
rlabel metal2 s 179758 -960 179870 480 8 la_data_in[15]
port 181 nsew signal input
rlabel metal2 s 183254 -960 183366 480 8 la_data_in[16]
port 182 nsew signal input
rlabel metal2 s 186842 -960 186954 480 8 la_data_in[17]
port 183 nsew signal input
rlabel metal2 s 190430 -960 190542 480 8 la_data_in[18]
port 184 nsew signal input
rlabel metal2 s 194018 -960 194130 480 8 la_data_in[19]
port 185 nsew signal input
rlabel metal2 s 129894 -960 130006 480 8 la_data_in[1]
port 186 nsew signal input
rlabel metal2 s 197514 -960 197626 480 8 la_data_in[20]
port 187 nsew signal input
rlabel metal2 s 201102 -960 201214 480 8 la_data_in[21]
port 188 nsew signal input
rlabel metal2 s 204690 -960 204802 480 8 la_data_in[22]
port 189 nsew signal input
rlabel metal2 s 208186 -960 208298 480 8 la_data_in[23]
port 190 nsew signal input
rlabel metal2 s 211774 -960 211886 480 8 la_data_in[24]
port 191 nsew signal input
rlabel metal2 s 215362 -960 215474 480 8 la_data_in[25]
port 192 nsew signal input
rlabel metal2 s 218950 -960 219062 480 8 la_data_in[26]
port 193 nsew signal input
rlabel metal2 s 222446 -960 222558 480 8 la_data_in[27]
port 194 nsew signal input
rlabel metal2 s 226034 -960 226146 480 8 la_data_in[28]
port 195 nsew signal input
rlabel metal2 s 229622 -960 229734 480 8 la_data_in[29]
port 196 nsew signal input
rlabel metal2 s 133482 -960 133594 480 8 la_data_in[2]
port 197 nsew signal input
rlabel metal2 s 233118 -960 233230 480 8 la_data_in[30]
port 198 nsew signal input
rlabel metal2 s 236706 -960 236818 480 8 la_data_in[31]
port 199 nsew signal input
rlabel metal2 s 240294 -960 240406 480 8 la_data_in[32]
port 200 nsew signal input
rlabel metal2 s 243882 -960 243994 480 8 la_data_in[33]
port 201 nsew signal input
rlabel metal2 s 247378 -960 247490 480 8 la_data_in[34]
port 202 nsew signal input
rlabel metal2 s 250966 -960 251078 480 8 la_data_in[35]
port 203 nsew signal input
rlabel metal2 s 254554 -960 254666 480 8 la_data_in[36]
port 204 nsew signal input
rlabel metal2 s 258050 -960 258162 480 8 la_data_in[37]
port 205 nsew signal input
rlabel metal2 s 261638 -960 261750 480 8 la_data_in[38]
port 206 nsew signal input
rlabel metal2 s 265226 -960 265338 480 8 la_data_in[39]
port 207 nsew signal input
rlabel metal2 s 136978 -960 137090 480 8 la_data_in[3]
port 208 nsew signal input
rlabel metal2 s 268722 -960 268834 480 8 la_data_in[40]
port 209 nsew signal input
rlabel metal2 s 272310 -960 272422 480 8 la_data_in[41]
port 210 nsew signal input
rlabel metal2 s 275898 -960 276010 480 8 la_data_in[42]
port 211 nsew signal input
rlabel metal2 s 279486 -960 279598 480 8 la_data_in[43]
port 212 nsew signal input
rlabel metal2 s 282982 -960 283094 480 8 la_data_in[44]
port 213 nsew signal input
rlabel metal2 s 286570 -960 286682 480 8 la_data_in[45]
port 214 nsew signal input
rlabel metal2 s 290158 -960 290270 480 8 la_data_in[46]
port 215 nsew signal input
rlabel metal2 s 293654 -960 293766 480 8 la_data_in[47]
port 216 nsew signal input
rlabel metal2 s 297242 -960 297354 480 8 la_data_in[48]
port 217 nsew signal input
rlabel metal2 s 300830 -960 300942 480 8 la_data_in[49]
port 218 nsew signal input
rlabel metal2 s 140566 -960 140678 480 8 la_data_in[4]
port 219 nsew signal input
rlabel metal2 s 304418 -960 304530 480 8 la_data_in[50]
port 220 nsew signal input
rlabel metal2 s 307914 -960 308026 480 8 la_data_in[51]
port 221 nsew signal input
rlabel metal2 s 311502 -960 311614 480 8 la_data_in[52]
port 222 nsew signal input
rlabel metal2 s 315090 -960 315202 480 8 la_data_in[53]
port 223 nsew signal input
rlabel metal2 s 318586 -960 318698 480 8 la_data_in[54]
port 224 nsew signal input
rlabel metal2 s 322174 -960 322286 480 8 la_data_in[55]
port 225 nsew signal input
rlabel metal2 s 325762 -960 325874 480 8 la_data_in[56]
port 226 nsew signal input
rlabel metal2 s 329258 -960 329370 480 8 la_data_in[57]
port 227 nsew signal input
rlabel metal2 s 332846 -960 332958 480 8 la_data_in[58]
port 228 nsew signal input
rlabel metal2 s 336434 -960 336546 480 8 la_data_in[59]
port 229 nsew signal input
rlabel metal2 s 144154 -960 144266 480 8 la_data_in[5]
port 230 nsew signal input
rlabel metal2 s 340022 -960 340134 480 8 la_data_in[60]
port 231 nsew signal input
rlabel metal2 s 343518 -960 343630 480 8 la_data_in[61]
port 232 nsew signal input
rlabel metal2 s 347106 -960 347218 480 8 la_data_in[62]
port 233 nsew signal input
rlabel metal2 s 350694 -960 350806 480 8 la_data_in[63]
port 234 nsew signal input
rlabel metal2 s 354190 -960 354302 480 8 la_data_in[64]
port 235 nsew signal input
rlabel metal2 s 357778 -960 357890 480 8 la_data_in[65]
port 236 nsew signal input
rlabel metal2 s 361366 -960 361478 480 8 la_data_in[66]
port 237 nsew signal input
rlabel metal2 s 364954 -960 365066 480 8 la_data_in[67]
port 238 nsew signal input
rlabel metal2 s 368450 -960 368562 480 8 la_data_in[68]
port 239 nsew signal input
rlabel metal2 s 372038 -960 372150 480 8 la_data_in[69]
port 240 nsew signal input
rlabel metal2 s 147650 -960 147762 480 8 la_data_in[6]
port 241 nsew signal input
rlabel metal2 s 375626 -960 375738 480 8 la_data_in[70]
port 242 nsew signal input
rlabel metal2 s 379122 -960 379234 480 8 la_data_in[71]
port 243 nsew signal input
rlabel metal2 s 382710 -960 382822 480 8 la_data_in[72]
port 244 nsew signal input
rlabel metal2 s 386298 -960 386410 480 8 la_data_in[73]
port 245 nsew signal input
rlabel metal2 s 389886 -960 389998 480 8 la_data_in[74]
port 246 nsew signal input
rlabel metal2 s 393382 -960 393494 480 8 la_data_in[75]
port 247 nsew signal input
rlabel metal2 s 396970 -960 397082 480 8 la_data_in[76]
port 248 nsew signal input
rlabel metal2 s 400558 -960 400670 480 8 la_data_in[77]
port 249 nsew signal input
rlabel metal2 s 404054 -960 404166 480 8 la_data_in[78]
port 250 nsew signal input
rlabel metal2 s 407642 -960 407754 480 8 la_data_in[79]
port 251 nsew signal input
rlabel metal2 s 151238 -960 151350 480 8 la_data_in[7]
port 252 nsew signal input
rlabel metal2 s 411230 -960 411342 480 8 la_data_in[80]
port 253 nsew signal input
rlabel metal2 s 414726 -960 414838 480 8 la_data_in[81]
port 254 nsew signal input
rlabel metal2 s 418314 -960 418426 480 8 la_data_in[82]
port 255 nsew signal input
rlabel metal2 s 421902 -960 422014 480 8 la_data_in[83]
port 256 nsew signal input
rlabel metal2 s 425490 -960 425602 480 8 la_data_in[84]
port 257 nsew signal input
rlabel metal2 s 428986 -960 429098 480 8 la_data_in[85]
port 258 nsew signal input
rlabel metal2 s 432574 -960 432686 480 8 la_data_in[86]
port 259 nsew signal input
rlabel metal2 s 436162 -960 436274 480 8 la_data_in[87]
port 260 nsew signal input
rlabel metal2 s 439658 -960 439770 480 8 la_data_in[88]
port 261 nsew signal input
rlabel metal2 s 443246 -960 443358 480 8 la_data_in[89]
port 262 nsew signal input
rlabel metal2 s 154826 -960 154938 480 8 la_data_in[8]
port 263 nsew signal input
rlabel metal2 s 446834 -960 446946 480 8 la_data_in[90]
port 264 nsew signal input
rlabel metal2 s 450422 -960 450534 480 8 la_data_in[91]
port 265 nsew signal input
rlabel metal2 s 453918 -960 454030 480 8 la_data_in[92]
port 266 nsew signal input
rlabel metal2 s 457506 -960 457618 480 8 la_data_in[93]
port 267 nsew signal input
rlabel metal2 s 461094 -960 461206 480 8 la_data_in[94]
port 268 nsew signal input
rlabel metal2 s 464590 -960 464702 480 8 la_data_in[95]
port 269 nsew signal input
rlabel metal2 s 468178 -960 468290 480 8 la_data_in[96]
port 270 nsew signal input
rlabel metal2 s 471766 -960 471878 480 8 la_data_in[97]
port 271 nsew signal input
rlabel metal2 s 475262 -960 475374 480 8 la_data_in[98]
port 272 nsew signal input
rlabel metal2 s 478850 -960 478962 480 8 la_data_in[99]
port 273 nsew signal input
rlabel metal2 s 158414 -960 158526 480 8 la_data_in[9]
port 274 nsew signal input
rlabel metal2 s 127502 -960 127614 480 8 la_data_out[0]
port 275 nsew signal output
rlabel metal2 s 483634 -960 483746 480 8 la_data_out[100]
port 276 nsew signal output
rlabel metal2 s 487222 -960 487334 480 8 la_data_out[101]
port 277 nsew signal output
rlabel metal2 s 490718 -960 490830 480 8 la_data_out[102]
port 278 nsew signal output
rlabel metal2 s 494306 -960 494418 480 8 la_data_out[103]
port 279 nsew signal output
rlabel metal2 s 497894 -960 498006 480 8 la_data_out[104]
port 280 nsew signal output
rlabel metal2 s 501390 -960 501502 480 8 la_data_out[105]
port 281 nsew signal output
rlabel metal2 s 504978 -960 505090 480 8 la_data_out[106]
port 282 nsew signal output
rlabel metal2 s 508566 -960 508678 480 8 la_data_out[107]
port 283 nsew signal output
rlabel metal2 s 512062 -960 512174 480 8 la_data_out[108]
port 284 nsew signal output
rlabel metal2 s 515650 -960 515762 480 8 la_data_out[109]
port 285 nsew signal output
rlabel metal2 s 163106 -960 163218 480 8 la_data_out[10]
port 286 nsew signal output
rlabel metal2 s 519238 -960 519350 480 8 la_data_out[110]
port 287 nsew signal output
rlabel metal2 s 522826 -960 522938 480 8 la_data_out[111]
port 288 nsew signal output
rlabel metal2 s 526322 -960 526434 480 8 la_data_out[112]
port 289 nsew signal output
rlabel metal2 s 529910 -960 530022 480 8 la_data_out[113]
port 290 nsew signal output
rlabel metal2 s 533498 -960 533610 480 8 la_data_out[114]
port 291 nsew signal output
rlabel metal2 s 536994 -960 537106 480 8 la_data_out[115]
port 292 nsew signal output
rlabel metal2 s 540582 -960 540694 480 8 la_data_out[116]
port 293 nsew signal output
rlabel metal2 s 544170 -960 544282 480 8 la_data_out[117]
port 294 nsew signal output
rlabel metal2 s 547758 -960 547870 480 8 la_data_out[118]
port 295 nsew signal output
rlabel metal2 s 551254 -960 551366 480 8 la_data_out[119]
port 296 nsew signal output
rlabel metal2 s 166694 -960 166806 480 8 la_data_out[11]
port 297 nsew signal output
rlabel metal2 s 554842 -960 554954 480 8 la_data_out[120]
port 298 nsew signal output
rlabel metal2 s 558430 -960 558542 480 8 la_data_out[121]
port 299 nsew signal output
rlabel metal2 s 561926 -960 562038 480 8 la_data_out[122]
port 300 nsew signal output
rlabel metal2 s 565514 -960 565626 480 8 la_data_out[123]
port 301 nsew signal output
rlabel metal2 s 569102 -960 569214 480 8 la_data_out[124]
port 302 nsew signal output
rlabel metal2 s 572598 -960 572710 480 8 la_data_out[125]
port 303 nsew signal output
rlabel metal2 s 576186 -960 576298 480 8 la_data_out[126]
port 304 nsew signal output
rlabel metal2 s 579774 -960 579886 480 8 la_data_out[127]
port 305 nsew signal output
rlabel metal2 s 170282 -960 170394 480 8 la_data_out[12]
port 306 nsew signal output
rlabel metal2 s 173778 -960 173890 480 8 la_data_out[13]
port 307 nsew signal output
rlabel metal2 s 177366 -960 177478 480 8 la_data_out[14]
port 308 nsew signal output
rlabel metal2 s 180954 -960 181066 480 8 la_data_out[15]
port 309 nsew signal output
rlabel metal2 s 184450 -960 184562 480 8 la_data_out[16]
port 310 nsew signal output
rlabel metal2 s 188038 -960 188150 480 8 la_data_out[17]
port 311 nsew signal output
rlabel metal2 s 191626 -960 191738 480 8 la_data_out[18]
port 312 nsew signal output
rlabel metal2 s 195214 -960 195326 480 8 la_data_out[19]
port 313 nsew signal output
rlabel metal2 s 131090 -960 131202 480 8 la_data_out[1]
port 314 nsew signal output
rlabel metal2 s 198710 -960 198822 480 8 la_data_out[20]
port 315 nsew signal output
rlabel metal2 s 202298 -960 202410 480 8 la_data_out[21]
port 316 nsew signal output
rlabel metal2 s 205886 -960 205998 480 8 la_data_out[22]
port 317 nsew signal output
rlabel metal2 s 209382 -960 209494 480 8 la_data_out[23]
port 318 nsew signal output
rlabel metal2 s 212970 -960 213082 480 8 la_data_out[24]
port 319 nsew signal output
rlabel metal2 s 216558 -960 216670 480 8 la_data_out[25]
port 320 nsew signal output
rlabel metal2 s 220054 -960 220166 480 8 la_data_out[26]
port 321 nsew signal output
rlabel metal2 s 223642 -960 223754 480 8 la_data_out[27]
port 322 nsew signal output
rlabel metal2 s 227230 -960 227342 480 8 la_data_out[28]
port 323 nsew signal output
rlabel metal2 s 230818 -960 230930 480 8 la_data_out[29]
port 324 nsew signal output
rlabel metal2 s 134586 -960 134698 480 8 la_data_out[2]
port 325 nsew signal output
rlabel metal2 s 234314 -960 234426 480 8 la_data_out[30]
port 326 nsew signal output
rlabel metal2 s 237902 -960 238014 480 8 la_data_out[31]
port 327 nsew signal output
rlabel metal2 s 241490 -960 241602 480 8 la_data_out[32]
port 328 nsew signal output
rlabel metal2 s 244986 -960 245098 480 8 la_data_out[33]
port 329 nsew signal output
rlabel metal2 s 248574 -960 248686 480 8 la_data_out[34]
port 330 nsew signal output
rlabel metal2 s 252162 -960 252274 480 8 la_data_out[35]
port 331 nsew signal output
rlabel metal2 s 255750 -960 255862 480 8 la_data_out[36]
port 332 nsew signal output
rlabel metal2 s 259246 -960 259358 480 8 la_data_out[37]
port 333 nsew signal output
rlabel metal2 s 262834 -960 262946 480 8 la_data_out[38]
port 334 nsew signal output
rlabel metal2 s 266422 -960 266534 480 8 la_data_out[39]
port 335 nsew signal output
rlabel metal2 s 138174 -960 138286 480 8 la_data_out[3]
port 336 nsew signal output
rlabel metal2 s 269918 -960 270030 480 8 la_data_out[40]
port 337 nsew signal output
rlabel metal2 s 273506 -960 273618 480 8 la_data_out[41]
port 338 nsew signal output
rlabel metal2 s 277094 -960 277206 480 8 la_data_out[42]
port 339 nsew signal output
rlabel metal2 s 280590 -960 280702 480 8 la_data_out[43]
port 340 nsew signal output
rlabel metal2 s 284178 -960 284290 480 8 la_data_out[44]
port 341 nsew signal output
rlabel metal2 s 287766 -960 287878 480 8 la_data_out[45]
port 342 nsew signal output
rlabel metal2 s 291354 -960 291466 480 8 la_data_out[46]
port 343 nsew signal output
rlabel metal2 s 294850 -960 294962 480 8 la_data_out[47]
port 344 nsew signal output
rlabel metal2 s 298438 -960 298550 480 8 la_data_out[48]
port 345 nsew signal output
rlabel metal2 s 302026 -960 302138 480 8 la_data_out[49]
port 346 nsew signal output
rlabel metal2 s 141762 -960 141874 480 8 la_data_out[4]
port 347 nsew signal output
rlabel metal2 s 305522 -960 305634 480 8 la_data_out[50]
port 348 nsew signal output
rlabel metal2 s 309110 -960 309222 480 8 la_data_out[51]
port 349 nsew signal output
rlabel metal2 s 312698 -960 312810 480 8 la_data_out[52]
port 350 nsew signal output
rlabel metal2 s 316286 -960 316398 480 8 la_data_out[53]
port 351 nsew signal output
rlabel metal2 s 319782 -960 319894 480 8 la_data_out[54]
port 352 nsew signal output
rlabel metal2 s 323370 -960 323482 480 8 la_data_out[55]
port 353 nsew signal output
rlabel metal2 s 326958 -960 327070 480 8 la_data_out[56]
port 354 nsew signal output
rlabel metal2 s 330454 -960 330566 480 8 la_data_out[57]
port 355 nsew signal output
rlabel metal2 s 334042 -960 334154 480 8 la_data_out[58]
port 356 nsew signal output
rlabel metal2 s 337630 -960 337742 480 8 la_data_out[59]
port 357 nsew signal output
rlabel metal2 s 145350 -960 145462 480 8 la_data_out[5]
port 358 nsew signal output
rlabel metal2 s 341218 -960 341330 480 8 la_data_out[60]
port 359 nsew signal output
rlabel metal2 s 344714 -960 344826 480 8 la_data_out[61]
port 360 nsew signal output
rlabel metal2 s 348302 -960 348414 480 8 la_data_out[62]
port 361 nsew signal output
rlabel metal2 s 351890 -960 352002 480 8 la_data_out[63]
port 362 nsew signal output
rlabel metal2 s 355386 -960 355498 480 8 la_data_out[64]
port 363 nsew signal output
rlabel metal2 s 358974 -960 359086 480 8 la_data_out[65]
port 364 nsew signal output
rlabel metal2 s 362562 -960 362674 480 8 la_data_out[66]
port 365 nsew signal output
rlabel metal2 s 366058 -960 366170 480 8 la_data_out[67]
port 366 nsew signal output
rlabel metal2 s 369646 -960 369758 480 8 la_data_out[68]
port 367 nsew signal output
rlabel metal2 s 373234 -960 373346 480 8 la_data_out[69]
port 368 nsew signal output
rlabel metal2 s 148846 -960 148958 480 8 la_data_out[6]
port 369 nsew signal output
rlabel metal2 s 376822 -960 376934 480 8 la_data_out[70]
port 370 nsew signal output
rlabel metal2 s 380318 -960 380430 480 8 la_data_out[71]
port 371 nsew signal output
rlabel metal2 s 383906 -960 384018 480 8 la_data_out[72]
port 372 nsew signal output
rlabel metal2 s 387494 -960 387606 480 8 la_data_out[73]
port 373 nsew signal output
rlabel metal2 s 390990 -960 391102 480 8 la_data_out[74]
port 374 nsew signal output
rlabel metal2 s 394578 -960 394690 480 8 la_data_out[75]
port 375 nsew signal output
rlabel metal2 s 398166 -960 398278 480 8 la_data_out[76]
port 376 nsew signal output
rlabel metal2 s 401754 -960 401866 480 8 la_data_out[77]
port 377 nsew signal output
rlabel metal2 s 405250 -960 405362 480 8 la_data_out[78]
port 378 nsew signal output
rlabel metal2 s 408838 -960 408950 480 8 la_data_out[79]
port 379 nsew signal output
rlabel metal2 s 152434 -960 152546 480 8 la_data_out[7]
port 380 nsew signal output
rlabel metal2 s 412426 -960 412538 480 8 la_data_out[80]
port 381 nsew signal output
rlabel metal2 s 415922 -960 416034 480 8 la_data_out[81]
port 382 nsew signal output
rlabel metal2 s 419510 -960 419622 480 8 la_data_out[82]
port 383 nsew signal output
rlabel metal2 s 423098 -960 423210 480 8 la_data_out[83]
port 384 nsew signal output
rlabel metal2 s 426594 -960 426706 480 8 la_data_out[84]
port 385 nsew signal output
rlabel metal2 s 430182 -960 430294 480 8 la_data_out[85]
port 386 nsew signal output
rlabel metal2 s 433770 -960 433882 480 8 la_data_out[86]
port 387 nsew signal output
rlabel metal2 s 437358 -960 437470 480 8 la_data_out[87]
port 388 nsew signal output
rlabel metal2 s 440854 -960 440966 480 8 la_data_out[88]
port 389 nsew signal output
rlabel metal2 s 444442 -960 444554 480 8 la_data_out[89]
port 390 nsew signal output
rlabel metal2 s 156022 -960 156134 480 8 la_data_out[8]
port 391 nsew signal output
rlabel metal2 s 448030 -960 448142 480 8 la_data_out[90]
port 392 nsew signal output
rlabel metal2 s 451526 -960 451638 480 8 la_data_out[91]
port 393 nsew signal output
rlabel metal2 s 455114 -960 455226 480 8 la_data_out[92]
port 394 nsew signal output
rlabel metal2 s 458702 -960 458814 480 8 la_data_out[93]
port 395 nsew signal output
rlabel metal2 s 462290 -960 462402 480 8 la_data_out[94]
port 396 nsew signal output
rlabel metal2 s 465786 -960 465898 480 8 la_data_out[95]
port 397 nsew signal output
rlabel metal2 s 469374 -960 469486 480 8 la_data_out[96]
port 398 nsew signal output
rlabel metal2 s 472962 -960 473074 480 8 la_data_out[97]
port 399 nsew signal output
rlabel metal2 s 476458 -960 476570 480 8 la_data_out[98]
port 400 nsew signal output
rlabel metal2 s 480046 -960 480158 480 8 la_data_out[99]
port 401 nsew signal output
rlabel metal2 s 159518 -960 159630 480 8 la_data_out[9]
port 402 nsew signal output
rlabel metal2 s 128698 -960 128810 480 8 la_oenb[0]
port 403 nsew signal input
rlabel metal2 s 484830 -960 484942 480 8 la_oenb[100]
port 404 nsew signal input
rlabel metal2 s 488326 -960 488438 480 8 la_oenb[101]
port 405 nsew signal input
rlabel metal2 s 491914 -960 492026 480 8 la_oenb[102]
port 406 nsew signal input
rlabel metal2 s 495502 -960 495614 480 8 la_oenb[103]
port 407 nsew signal input
rlabel metal2 s 499090 -960 499202 480 8 la_oenb[104]
port 408 nsew signal input
rlabel metal2 s 502586 -960 502698 480 8 la_oenb[105]
port 409 nsew signal input
rlabel metal2 s 506174 -960 506286 480 8 la_oenb[106]
port 410 nsew signal input
rlabel metal2 s 509762 -960 509874 480 8 la_oenb[107]
port 411 nsew signal input
rlabel metal2 s 513258 -960 513370 480 8 la_oenb[108]
port 412 nsew signal input
rlabel metal2 s 516846 -960 516958 480 8 la_oenb[109]
port 413 nsew signal input
rlabel metal2 s 164302 -960 164414 480 8 la_oenb[10]
port 414 nsew signal input
rlabel metal2 s 520434 -960 520546 480 8 la_oenb[110]
port 415 nsew signal input
rlabel metal2 s 523930 -960 524042 480 8 la_oenb[111]
port 416 nsew signal input
rlabel metal2 s 527518 -960 527630 480 8 la_oenb[112]
port 417 nsew signal input
rlabel metal2 s 531106 -960 531218 480 8 la_oenb[113]
port 418 nsew signal input
rlabel metal2 s 534694 -960 534806 480 8 la_oenb[114]
port 419 nsew signal input
rlabel metal2 s 538190 -960 538302 480 8 la_oenb[115]
port 420 nsew signal input
rlabel metal2 s 541778 -960 541890 480 8 la_oenb[116]
port 421 nsew signal input
rlabel metal2 s 545366 -960 545478 480 8 la_oenb[117]
port 422 nsew signal input
rlabel metal2 s 548862 -960 548974 480 8 la_oenb[118]
port 423 nsew signal input
rlabel metal2 s 552450 -960 552562 480 8 la_oenb[119]
port 424 nsew signal input
rlabel metal2 s 167890 -960 168002 480 8 la_oenb[11]
port 425 nsew signal input
rlabel metal2 s 556038 -960 556150 480 8 la_oenb[120]
port 426 nsew signal input
rlabel metal2 s 559626 -960 559738 480 8 la_oenb[121]
port 427 nsew signal input
rlabel metal2 s 563122 -960 563234 480 8 la_oenb[122]
port 428 nsew signal input
rlabel metal2 s 566710 -960 566822 480 8 la_oenb[123]
port 429 nsew signal input
rlabel metal2 s 570298 -960 570410 480 8 la_oenb[124]
port 430 nsew signal input
rlabel metal2 s 573794 -960 573906 480 8 la_oenb[125]
port 431 nsew signal input
rlabel metal2 s 577382 -960 577494 480 8 la_oenb[126]
port 432 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 la_oenb[127]
port 433 nsew signal input
rlabel metal2 s 171386 -960 171498 480 8 la_oenb[12]
port 434 nsew signal input
rlabel metal2 s 174974 -960 175086 480 8 la_oenb[13]
port 435 nsew signal input
rlabel metal2 s 178562 -960 178674 480 8 la_oenb[14]
port 436 nsew signal input
rlabel metal2 s 182150 -960 182262 480 8 la_oenb[15]
port 437 nsew signal input
rlabel metal2 s 185646 -960 185758 480 8 la_oenb[16]
port 438 nsew signal input
rlabel metal2 s 189234 -960 189346 480 8 la_oenb[17]
port 439 nsew signal input
rlabel metal2 s 192822 -960 192934 480 8 la_oenb[18]
port 440 nsew signal input
rlabel metal2 s 196318 -960 196430 480 8 la_oenb[19]
port 441 nsew signal input
rlabel metal2 s 132286 -960 132398 480 8 la_oenb[1]
port 442 nsew signal input
rlabel metal2 s 199906 -960 200018 480 8 la_oenb[20]
port 443 nsew signal input
rlabel metal2 s 203494 -960 203606 480 8 la_oenb[21]
port 444 nsew signal input
rlabel metal2 s 207082 -960 207194 480 8 la_oenb[22]
port 445 nsew signal input
rlabel metal2 s 210578 -960 210690 480 8 la_oenb[23]
port 446 nsew signal input
rlabel metal2 s 214166 -960 214278 480 8 la_oenb[24]
port 447 nsew signal input
rlabel metal2 s 217754 -960 217866 480 8 la_oenb[25]
port 448 nsew signal input
rlabel metal2 s 221250 -960 221362 480 8 la_oenb[26]
port 449 nsew signal input
rlabel metal2 s 224838 -960 224950 480 8 la_oenb[27]
port 450 nsew signal input
rlabel metal2 s 228426 -960 228538 480 8 la_oenb[28]
port 451 nsew signal input
rlabel metal2 s 231922 -960 232034 480 8 la_oenb[29]
port 452 nsew signal input
rlabel metal2 s 135782 -960 135894 480 8 la_oenb[2]
port 453 nsew signal input
rlabel metal2 s 235510 -960 235622 480 8 la_oenb[30]
port 454 nsew signal input
rlabel metal2 s 239098 -960 239210 480 8 la_oenb[31]
port 455 nsew signal input
rlabel metal2 s 242686 -960 242798 480 8 la_oenb[32]
port 456 nsew signal input
rlabel metal2 s 246182 -960 246294 480 8 la_oenb[33]
port 457 nsew signal input
rlabel metal2 s 249770 -960 249882 480 8 la_oenb[34]
port 458 nsew signal input
rlabel metal2 s 253358 -960 253470 480 8 la_oenb[35]
port 459 nsew signal input
rlabel metal2 s 256854 -960 256966 480 8 la_oenb[36]
port 460 nsew signal input
rlabel metal2 s 260442 -960 260554 480 8 la_oenb[37]
port 461 nsew signal input
rlabel metal2 s 264030 -960 264142 480 8 la_oenb[38]
port 462 nsew signal input
rlabel metal2 s 267618 -960 267730 480 8 la_oenb[39]
port 463 nsew signal input
rlabel metal2 s 139370 -960 139482 480 8 la_oenb[3]
port 464 nsew signal input
rlabel metal2 s 271114 -960 271226 480 8 la_oenb[40]
port 465 nsew signal input
rlabel metal2 s 274702 -960 274814 480 8 la_oenb[41]
port 466 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_oenb[42]
port 467 nsew signal input
rlabel metal2 s 281786 -960 281898 480 8 la_oenb[43]
port 468 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_oenb[44]
port 469 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_oenb[45]
port 470 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_oenb[46]
port 471 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_oenb[47]
port 472 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_oenb[48]
port 473 nsew signal input
rlabel metal2 s 303222 -960 303334 480 8 la_oenb[49]
port 474 nsew signal input
rlabel metal2 s 142958 -960 143070 480 8 la_oenb[4]
port 475 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_oenb[50]
port 476 nsew signal input
rlabel metal2 s 310306 -960 310418 480 8 la_oenb[51]
port 477 nsew signal input
rlabel metal2 s 313894 -960 314006 480 8 la_oenb[52]
port 478 nsew signal input
rlabel metal2 s 317390 -960 317502 480 8 la_oenb[53]
port 479 nsew signal input
rlabel metal2 s 320978 -960 321090 480 8 la_oenb[54]
port 480 nsew signal input
rlabel metal2 s 324566 -960 324678 480 8 la_oenb[55]
port 481 nsew signal input
rlabel metal2 s 328154 -960 328266 480 8 la_oenb[56]
port 482 nsew signal input
rlabel metal2 s 331650 -960 331762 480 8 la_oenb[57]
port 483 nsew signal input
rlabel metal2 s 335238 -960 335350 480 8 la_oenb[58]
port 484 nsew signal input
rlabel metal2 s 338826 -960 338938 480 8 la_oenb[59]
port 485 nsew signal input
rlabel metal2 s 146546 -960 146658 480 8 la_oenb[5]
port 486 nsew signal input
rlabel metal2 s 342322 -960 342434 480 8 la_oenb[60]
port 487 nsew signal input
rlabel metal2 s 345910 -960 346022 480 8 la_oenb[61]
port 488 nsew signal input
rlabel metal2 s 349498 -960 349610 480 8 la_oenb[62]
port 489 nsew signal input
rlabel metal2 s 353086 -960 353198 480 8 la_oenb[63]
port 490 nsew signal input
rlabel metal2 s 356582 -960 356694 480 8 la_oenb[64]
port 491 nsew signal input
rlabel metal2 s 360170 -960 360282 480 8 la_oenb[65]
port 492 nsew signal input
rlabel metal2 s 363758 -960 363870 480 8 la_oenb[66]
port 493 nsew signal input
rlabel metal2 s 367254 -960 367366 480 8 la_oenb[67]
port 494 nsew signal input
rlabel metal2 s 370842 -960 370954 480 8 la_oenb[68]
port 495 nsew signal input
rlabel metal2 s 374430 -960 374542 480 8 la_oenb[69]
port 496 nsew signal input
rlabel metal2 s 150042 -960 150154 480 8 la_oenb[6]
port 497 nsew signal input
rlabel metal2 s 377926 -960 378038 480 8 la_oenb[70]
port 498 nsew signal input
rlabel metal2 s 381514 -960 381626 480 8 la_oenb[71]
port 499 nsew signal input
rlabel metal2 s 385102 -960 385214 480 8 la_oenb[72]
port 500 nsew signal input
rlabel metal2 s 388690 -960 388802 480 8 la_oenb[73]
port 501 nsew signal input
rlabel metal2 s 392186 -960 392298 480 8 la_oenb[74]
port 502 nsew signal input
rlabel metal2 s 395774 -960 395886 480 8 la_oenb[75]
port 503 nsew signal input
rlabel metal2 s 399362 -960 399474 480 8 la_oenb[76]
port 504 nsew signal input
rlabel metal2 s 402858 -960 402970 480 8 la_oenb[77]
port 505 nsew signal input
rlabel metal2 s 406446 -960 406558 480 8 la_oenb[78]
port 506 nsew signal input
rlabel metal2 s 410034 -960 410146 480 8 la_oenb[79]
port 507 nsew signal input
rlabel metal2 s 153630 -960 153742 480 8 la_oenb[7]
port 508 nsew signal input
rlabel metal2 s 413622 -960 413734 480 8 la_oenb[80]
port 509 nsew signal input
rlabel metal2 s 417118 -960 417230 480 8 la_oenb[81]
port 510 nsew signal input
rlabel metal2 s 420706 -960 420818 480 8 la_oenb[82]
port 511 nsew signal input
rlabel metal2 s 424294 -960 424406 480 8 la_oenb[83]
port 512 nsew signal input
rlabel metal2 s 427790 -960 427902 480 8 la_oenb[84]
port 513 nsew signal input
rlabel metal2 s 431378 -960 431490 480 8 la_oenb[85]
port 514 nsew signal input
rlabel metal2 s 434966 -960 435078 480 8 la_oenb[86]
port 515 nsew signal input
rlabel metal2 s 438554 -960 438666 480 8 la_oenb[87]
port 516 nsew signal input
rlabel metal2 s 442050 -960 442162 480 8 la_oenb[88]
port 517 nsew signal input
rlabel metal2 s 445638 -960 445750 480 8 la_oenb[89]
port 518 nsew signal input
rlabel metal2 s 157218 -960 157330 480 8 la_oenb[8]
port 519 nsew signal input
rlabel metal2 s 449226 -960 449338 480 8 la_oenb[90]
port 520 nsew signal input
rlabel metal2 s 452722 -960 452834 480 8 la_oenb[91]
port 521 nsew signal input
rlabel metal2 s 456310 -960 456422 480 8 la_oenb[92]
port 522 nsew signal input
rlabel metal2 s 459898 -960 460010 480 8 la_oenb[93]
port 523 nsew signal input
rlabel metal2 s 463394 -960 463506 480 8 la_oenb[94]
port 524 nsew signal input
rlabel metal2 s 466982 -960 467094 480 8 la_oenb[95]
port 525 nsew signal input
rlabel metal2 s 470570 -960 470682 480 8 la_oenb[96]
port 526 nsew signal input
rlabel metal2 s 474158 -960 474270 480 8 la_oenb[97]
port 527 nsew signal input
rlabel metal2 s 477654 -960 477766 480 8 la_oenb[98]
port 528 nsew signal input
rlabel metal2 s 481242 -960 481354 480 8 la_oenb[99]
port 529 nsew signal input
rlabel metal2 s 160714 -960 160826 480 8 la_oenb[9]
port 530 nsew signal input
rlabel metal2 s 582166 -960 582278 480 8 user_clock2
port 531 nsew signal input
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 -1894 218414 198000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 -1894 254414 198000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 -1894 290414 198000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 -1894 326414 198000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 -1894 362414 198000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 322000 218414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 322000 254414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 322000 290414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 322000 326414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 322000 362414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 533 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 -3814 222134 198000 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 -3814 258134 198000 6 vccd2
port 533 nsew power input
rlabel metal4 s 293514 -3814 294134 198000 6 vccd2
port 533 nsew power input
rlabel metal4 s 329514 -3814 330134 198000 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 -3814 366134 198000 6 vccd2
port 533 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 322000 222134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 322000 258134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 293514 322000 294134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 329514 322000 330134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 322000 366134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 533 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 534 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 -5734 225854 198000 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 -5734 261854 198000 6 vdda1
port 534 nsew power input
rlabel metal4 s 297234 -5734 297854 198000 6 vdda1
port 534 nsew power input
rlabel metal4 s 333234 -5734 333854 198000 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 -5734 369854 198000 6 vdda1
port 534 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 322000 225854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 322000 261854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 297234 322000 297854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 333234 322000 333854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 322000 369854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 534 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 535 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 -7654 229574 198000 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 -7654 265574 198000 6 vdda2
port 535 nsew power input
rlabel metal4 s 300954 -7654 301574 198000 6 vdda2
port 535 nsew power input
rlabel metal4 s 336954 -7654 337574 198000 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 -7654 373574 198000 6 vdda2
port 535 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 322000 229574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 322000 265574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 300954 322000 301574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 336954 322000 337574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 322000 373574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 535 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 207234 -5734 207854 198000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 -5734 243854 198000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 -5734 279854 198000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 315234 -5734 315854 198000 6 vssa1
port 536 nsew ground input
rlabel metal4 s 351234 -5734 351854 198000 6 vssa1
port 536 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 207234 322000 207854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 322000 243854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 322000 279854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 315234 322000 315854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 351234 322000 351854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 210954 -7654 211574 198000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 -7654 247574 198000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 -7654 283574 198000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 318954 -7654 319574 198000 6 vssa2
port 537 nsew ground input
rlabel metal4 s 354954 -7654 355574 198000 6 vssa2
port 537 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 210954 322000 211574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 322000 247574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 322000 283574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 318954 322000 319574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 354954 322000 355574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 199794 -1894 200414 198000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 -1894 236414 198000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 -1894 272414 198000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 307794 -1894 308414 198000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 343794 -1894 344414 198000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 -1894 380414 198000 6 vssd1
port 538 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 199794 322000 200414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 322000 236414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 322000 272414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 307794 322000 308414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 343794 322000 344414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 322000 380414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 203514 -3814 204134 198000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 -3814 240134 198000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 -3814 276134 198000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 311514 -3814 312134 198000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 347514 -3814 348134 198000 6 vssd2
port 539 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 203514 322000 204134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 322000 240134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 322000 276134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 311514 322000 312134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 347514 322000 348134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 48014 -960 48126 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51510 -960 51622 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 55098 -960 55210 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58686 -960 58798 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 62182 -960 62294 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65770 -960 65882 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69358 -960 69470 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72946 -960 73058 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76442 -960 76554 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 80030 -960 80142 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83618 -960 83730 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 87114 -960 87226 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90702 -960 90814 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 94290 -960 94402 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97878 -960 97990 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101374 -960 101486 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104962 -960 105074 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108550 -960 108662 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 112046 -960 112158 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115634 -960 115746 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17102 -960 17214 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 119222 -960 119334 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122718 -960 122830 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26578 -960 26690 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30166 -960 30278 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33754 -960 33866 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37250 -960 37362 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40838 -960 40950 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44426 -960 44538 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 49210 -960 49322 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52706 -960 52818 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56294 -960 56406 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59882 -960 59994 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63378 -960 63490 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66966 -960 67078 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70554 -960 70666 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 74050 -960 74162 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77638 -960 77750 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 81226 -960 81338 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84814 -960 84926 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 88310 -960 88422 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91898 -960 92010 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95486 -960 95598 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98982 -960 99094 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102570 -960 102682 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 106158 -960 106270 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109746 -960 109858 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 113242 -960 113354 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116830 -960 116942 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 120418 -960 120530 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123914 -960 124026 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27774 -960 27886 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31362 -960 31474 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38446 -960 38558 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 42034 -960 42146 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45622 -960 45734 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50314 -960 50426 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53902 -960 54014 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57490 -960 57602 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 61078 -960 61190 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64574 -960 64686 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 68162 -960 68274 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71750 -960 71862 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 75246 -960 75358 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78834 -960 78946 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82422 -960 82534 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85918 -960 86030 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89506 -960 89618 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 93094 -960 93206 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96682 -960 96794 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 100178 -960 100290 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103766 -960 103878 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 107354 -960 107466 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110850 -960 110962 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 114438 -960 114550 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 118026 -960 118138 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121614 -960 121726 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 125110 -960 125222 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28970 -960 29082 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32558 -960 32670 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39642 -960 39754 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43230 -960 43342 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46818 -960 46930 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25382 -960 25494 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8510836
string GDS_FILE /opt/caravel/caravel_example/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 6778572
<< end >>

