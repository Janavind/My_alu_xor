VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 130.600 900.000 131.200 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 596.000 196.790 600.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 596.000 478.310 600.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 430.480 900.000 431.080 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 596.000 253.370 600.000 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 596.000 534.430 600.000 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 467.880 900.000 468.480 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END A1[7]
  PIN ALU_Out1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 55.800 900.000 56.400 ;
    END
  END ALU_Out1[0]
  PIN ALU_Out1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END ALU_Out1[1]
  PIN ALU_Out1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END ALU_Out1[2]
  PIN ALU_Out1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 280.200 900.000 280.800 ;
    END
  END ALU_Out1[3]
  PIN ALU_Out1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 355.680 900.000 356.280 ;
    END
  END ALU_Out1[4]
  PIN ALU_Out1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END ALU_Out1[5]
  PIN ALU_Out1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 509.360 4.000 509.960 ;
    END
  END ALU_Out1[6]
  PIN ALU_Out1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END ALU_Out1[7]
  PIN ALU_Out2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END ALU_Out2[0]
  PIN ALU_Out2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END ALU_Out2[1]
  PIN ALU_Out2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 205.400 900.000 206.000 ;
    END
  END ALU_Out2[2]
  PIN ALU_Out2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END ALU_Out2[3]
  PIN ALU_Out2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 596.000 591.010 600.000 ;
    END
  END ALU_Out2[4]
  PIN ALU_Out2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END ALU_Out2[5]
  PIN ALU_Out2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 596.000 815.950 600.000 ;
    END
  END ALU_Out2[6]
  PIN ALU_Out2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.200 4.000 569.800 ;
    END
  END ALU_Out2[7]
  PIN ALU_Sel1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END ALU_Sel1[0]
  PIN ALU_Sel1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END ALU_Sel1[1]
  PIN ALU_Sel2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 596.000 28.430 600.000 ;
    END
  END ALU_Sel2[0]
  PIN ALU_Sel2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 596.000 140.670 600.000 ;
    END
  END ALU_Sel2[1]
  PIN B0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 93.200 900.000 93.800 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 596.000 365.610 600.000 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 596.000 647.130 600.000 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 505.280 900.000 505.880 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 596.000 872.070 600.000 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 168.000 900.000 168.600 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 596.000 309.490 600.000 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 596.000 422.190 600.000 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 393.080 900.000 393.680 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 596.000 759.830 600.000 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 542.680 900.000 543.280 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END B1[7]
  PIN CarryOut1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END CarryOut1
  PIN CarryOut2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 18.400 900.000 19.000 ;
    END
  END CarryOut2
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END clk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 596.000 84.550 600.000 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 242.800 900.000 243.400 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 318.280 900.000 318.880 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 596.000 703.250 600.000 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 580.080 900.000 580.680 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END x[7]
  PIN y
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END y
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 8.540 894.240 587.760 ;
      LAYER met2 ;
        RECT 6.990 595.720 27.870 596.770 ;
        RECT 28.710 595.720 83.990 596.770 ;
        RECT 84.830 595.720 140.110 596.770 ;
        RECT 140.950 595.720 196.230 596.770 ;
        RECT 197.070 595.720 252.810 596.770 ;
        RECT 253.650 595.720 308.930 596.770 ;
        RECT 309.770 595.720 365.050 596.770 ;
        RECT 365.890 595.720 421.630 596.770 ;
        RECT 422.470 595.720 477.750 596.770 ;
        RECT 478.590 595.720 533.870 596.770 ;
        RECT 534.710 595.720 590.450 596.770 ;
        RECT 591.290 595.720 646.570 596.770 ;
        RECT 647.410 595.720 702.690 596.770 ;
        RECT 703.530 595.720 759.270 596.770 ;
        RECT 760.110 595.720 815.390 596.770 ;
        RECT 816.230 595.720 871.510 596.770 ;
        RECT 872.350 595.720 890.930 596.770 ;
        RECT 6.990 4.280 890.930 595.720 ;
        RECT 6.990 4.000 20.050 4.280 ;
        RECT 20.890 4.000 60.530 4.280 ;
        RECT 61.370 4.000 101.470 4.280 ;
        RECT 102.310 4.000 142.410 4.280 ;
        RECT 143.250 4.000 183.350 4.280 ;
        RECT 184.190 4.000 224.290 4.280 ;
        RECT 225.130 4.000 265.230 4.280 ;
        RECT 266.070 4.000 306.170 4.280 ;
        RECT 307.010 4.000 347.110 4.280 ;
        RECT 347.950 4.000 388.050 4.280 ;
        RECT 388.890 4.000 428.990 4.280 ;
        RECT 429.830 4.000 469.930 4.280 ;
        RECT 470.770 4.000 510.870 4.280 ;
        RECT 511.710 4.000 551.810 4.280 ;
        RECT 552.650 4.000 592.750 4.280 ;
        RECT 593.590 4.000 633.690 4.280 ;
        RECT 634.530 4.000 674.630 4.280 ;
        RECT 675.470 4.000 715.570 4.280 ;
        RECT 716.410 4.000 756.510 4.280 ;
        RECT 757.350 4.000 797.450 4.280 ;
        RECT 798.290 4.000 838.390 4.280 ;
        RECT 839.230 4.000 879.330 4.280 ;
        RECT 880.170 4.000 890.930 4.280 ;
      LAYER met3 ;
        RECT 4.000 581.080 896.000 587.685 ;
        RECT 4.000 579.680 895.600 581.080 ;
        RECT 4.000 570.200 896.000 579.680 ;
        RECT 4.400 568.800 896.000 570.200 ;
        RECT 4.000 543.680 896.000 568.800 ;
        RECT 4.000 542.280 895.600 543.680 ;
        RECT 4.000 510.360 896.000 542.280 ;
        RECT 4.400 508.960 896.000 510.360 ;
        RECT 4.000 506.280 896.000 508.960 ;
        RECT 4.000 504.880 895.600 506.280 ;
        RECT 4.000 468.880 896.000 504.880 ;
        RECT 4.000 467.480 895.600 468.880 ;
        RECT 4.000 450.520 896.000 467.480 ;
        RECT 4.400 449.120 896.000 450.520 ;
        RECT 4.000 431.480 896.000 449.120 ;
        RECT 4.000 430.080 895.600 431.480 ;
        RECT 4.000 394.080 896.000 430.080 ;
        RECT 4.000 392.680 895.600 394.080 ;
        RECT 4.000 390.680 896.000 392.680 ;
        RECT 4.400 389.280 896.000 390.680 ;
        RECT 4.000 356.680 896.000 389.280 ;
        RECT 4.000 355.280 895.600 356.680 ;
        RECT 4.000 330.840 896.000 355.280 ;
        RECT 4.400 329.440 896.000 330.840 ;
        RECT 4.000 319.280 896.000 329.440 ;
        RECT 4.000 317.880 895.600 319.280 ;
        RECT 4.000 281.200 896.000 317.880 ;
        RECT 4.000 279.800 895.600 281.200 ;
        RECT 4.000 270.320 896.000 279.800 ;
        RECT 4.400 268.920 896.000 270.320 ;
        RECT 4.000 243.800 896.000 268.920 ;
        RECT 4.000 242.400 895.600 243.800 ;
        RECT 4.000 210.480 896.000 242.400 ;
        RECT 4.400 209.080 896.000 210.480 ;
        RECT 4.000 206.400 896.000 209.080 ;
        RECT 4.000 205.000 895.600 206.400 ;
        RECT 4.000 169.000 896.000 205.000 ;
        RECT 4.000 167.600 895.600 169.000 ;
        RECT 4.000 150.640 896.000 167.600 ;
        RECT 4.400 149.240 896.000 150.640 ;
        RECT 4.000 131.600 896.000 149.240 ;
        RECT 4.000 130.200 895.600 131.600 ;
        RECT 4.000 94.200 896.000 130.200 ;
        RECT 4.000 92.800 895.600 94.200 ;
        RECT 4.000 90.800 896.000 92.800 ;
        RECT 4.400 89.400 896.000 90.800 ;
        RECT 4.000 56.800 896.000 89.400 ;
        RECT 4.000 55.400 895.600 56.800 ;
        RECT 4.000 30.960 896.000 55.400 ;
        RECT 4.400 29.560 896.000 30.960 ;
        RECT 4.000 19.400 896.000 29.560 ;
        RECT 4.000 18.000 895.600 19.400 ;
        RECT 4.000 10.715 896.000 18.000 ;
      LAYER met4 ;
        RECT 473.175 210.295 481.440 283.385 ;
        RECT 483.840 210.295 511.225 283.385 ;
  END
END user_proj_example
END LIBRARY

