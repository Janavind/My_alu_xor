magic
tech sky130A
magscale 1 2
timestamp 1647270986
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 1912 178848 117552
<< metal2 >>
rect 4250 119200 4306 120000
rect 12806 119200 12862 120000
rect 21362 119200 21418 120000
rect 29918 119200 29974 120000
rect 38474 119200 38530 120000
rect 47030 119200 47086 120000
rect 55678 119200 55734 120000
rect 64234 119200 64290 120000
rect 72790 119200 72846 120000
rect 81346 119200 81402 120000
rect 89902 119200 89958 120000
rect 98550 119200 98606 120000
rect 107106 119200 107162 120000
rect 115662 119200 115718 120000
rect 124218 119200 124274 120000
rect 132774 119200 132830 120000
rect 141422 119200 141478 120000
rect 149978 119200 150034 120000
rect 158534 119200 158590 120000
rect 167090 119200 167146 120000
rect 175646 119200 175702 120000
rect 4986 0 5042 800
rect 14922 0 14978 800
rect 24950 0 25006 800
rect 34978 0 35034 800
rect 44914 0 44970 800
rect 54942 0 54998 800
rect 64970 0 65026 800
rect 74998 0 75054 800
rect 84934 0 84990 800
rect 94962 0 95018 800
rect 104990 0 105046 800
rect 114926 0 114982 800
rect 124954 0 125010 800
rect 134982 0 135038 800
rect 145010 0 145066 800
rect 154946 0 155002 800
rect 164974 0 165030 800
rect 175002 0 175058 800
<< obsm2 >>
rect 1398 119144 4194 119354
rect 4362 119144 12750 119354
rect 12918 119144 21306 119354
rect 21474 119144 29862 119354
rect 30030 119144 38418 119354
rect 38586 119144 46974 119354
rect 47142 119144 55622 119354
rect 55790 119144 64178 119354
rect 64346 119144 72734 119354
rect 72902 119144 81290 119354
rect 81458 119144 89846 119354
rect 90014 119144 98494 119354
rect 98662 119144 107050 119354
rect 107218 119144 115606 119354
rect 115774 119144 124162 119354
rect 124330 119144 132718 119354
rect 132886 119144 141366 119354
rect 141534 119144 149922 119354
rect 150090 119144 158478 119354
rect 158646 119144 167034 119354
rect 167202 119144 175590 119354
rect 175758 119144 178186 119354
rect 1398 856 178186 119144
rect 1398 800 4930 856
rect 5098 800 14866 856
rect 15034 800 24894 856
rect 25062 800 34922 856
rect 35090 800 44858 856
rect 45026 800 54886 856
rect 55054 800 64914 856
rect 65082 800 74942 856
rect 75110 800 84878 856
rect 85046 800 94906 856
rect 95074 800 104934 856
rect 105102 800 114870 856
rect 115038 800 124898 856
rect 125066 800 134926 856
rect 135094 800 144954 856
rect 145122 800 154890 856
rect 155058 800 164918 856
rect 165086 800 174946 856
rect 175114 800 178186 856
<< metal3 >>
rect 179200 115608 180000 115728
rect 0 114384 800 114504
rect 179200 107040 180000 107160
rect 0 103504 800 103624
rect 179200 98472 180000 98592
rect 0 92624 800 92744
rect 179200 89904 180000 90024
rect 0 81744 800 81864
rect 179200 81336 180000 81456
rect 179200 72768 180000 72888
rect 0 70864 800 70984
rect 179200 64200 180000 64320
rect 0 59848 800 59968
rect 179200 55632 180000 55752
rect 0 48968 800 49088
rect 179200 47064 180000 47184
rect 179200 38496 180000 38616
rect 0 38088 800 38208
rect 179200 29928 180000 30048
rect 0 27208 800 27328
rect 179200 21360 180000 21480
rect 0 16328 800 16448
rect 179200 12792 180000 12912
rect 0 5448 800 5568
rect 179200 4224 180000 4344
<< obsm3 >>
rect 800 115808 179200 117537
rect 800 115528 179120 115808
rect 800 114584 179200 115528
rect 880 114304 179200 114584
rect 800 107240 179200 114304
rect 800 106960 179120 107240
rect 800 103704 179200 106960
rect 880 103424 179200 103704
rect 800 98672 179200 103424
rect 800 98392 179120 98672
rect 800 92824 179200 98392
rect 880 92544 179200 92824
rect 800 90104 179200 92544
rect 800 89824 179120 90104
rect 800 81944 179200 89824
rect 880 81664 179200 81944
rect 800 81536 179200 81664
rect 800 81256 179120 81536
rect 800 72968 179200 81256
rect 800 72688 179120 72968
rect 800 71064 179200 72688
rect 880 70784 179200 71064
rect 800 64400 179200 70784
rect 800 64120 179120 64400
rect 800 60048 179200 64120
rect 880 59768 179200 60048
rect 800 55832 179200 59768
rect 800 55552 179120 55832
rect 800 49168 179200 55552
rect 880 48888 179200 49168
rect 800 47264 179200 48888
rect 800 46984 179120 47264
rect 800 38696 179200 46984
rect 800 38416 179120 38696
rect 800 38288 179200 38416
rect 880 38008 179200 38288
rect 800 30128 179200 38008
rect 800 29848 179120 30128
rect 800 27408 179200 29848
rect 880 27128 179200 27408
rect 800 21560 179200 27128
rect 800 21280 179120 21560
rect 800 16528 179200 21280
rect 880 16248 179200 16528
rect 800 12992 179200 16248
rect 800 12712 179120 12992
rect 800 5648 179200 12712
rect 880 5368 179200 5648
rect 800 4424 179200 5368
rect 800 4144 179120 4424
rect 800 2143 179200 4144
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 89483 4659 96288 75309
rect 96768 4659 99669 75309
<< labels >>
rlabel metal2 s 14922 0 14978 800 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 179200 38496 180000 38616 6 A0[1]
port 2 nsew signal input
rlabel metal2 s 64234 119200 64290 120000 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 179200 72768 180000 72888 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 A0[4]
port 5 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 A0[5]
port 6 nsew signal input
rlabel metal2 s 149978 119200 150034 120000 6 A0[6]
port 7 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 A1[0]
port 9 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 A1[1]
port 10 nsew signal input
rlabel metal2 s 72790 119200 72846 120000 6 A1[2]
port 11 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 A1[3]
port 12 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 A1[4]
port 13 nsew signal input
rlabel metal2 s 115662 119200 115718 120000 6 A1[5]
port 14 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 A1[6]
port 15 nsew signal input
rlabel metal2 s 167090 119200 167146 120000 6 A1[7]
port 16 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 ALU_Out1[0]
port 17 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 ALU_Out1[1]
port 18 nsew signal output
rlabel metal3 s 179200 55632 180000 55752 6 ALU_Out1[2]
port 19 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 ALU_Out1[3]
port 20 nsew signal output
rlabel metal2 s 98550 119200 98606 120000 6 ALU_Out1[4]
port 21 nsew signal output
rlabel metal2 s 124218 119200 124274 120000 6 ALU_Out1[5]
port 22 nsew signal output
rlabel metal2 s 158534 119200 158590 120000 6 ALU_Out1[6]
port 23 nsew signal output
rlabel metal2 s 175646 119200 175702 120000 6 ALU_Out1[7]
port 24 nsew signal output
rlabel metal2 s 21362 119200 21418 120000 6 ALU_Out2[0]
port 25 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 ALU_Out2[1]
port 26 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 ALU_Out2[2]
port 27 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 ALU_Out2[3]
port 28 nsew signal output
rlabel metal3 s 179200 81336 180000 81456 6 ALU_Out2[4]
port 29 nsew signal output
rlabel metal3 s 0 81744 800 81864 6 ALU_Out2[5]
port 30 nsew signal output
rlabel metal3 s 179200 107040 180000 107160 6 ALU_Out2[6]
port 31 nsew signal output
rlabel metal3 s 179200 115608 180000 115728 6 ALU_Out2[7]
port 32 nsew signal output
rlabel metal3 s 179200 12792 180000 12912 6 ALU_Sel1[0]
port 33 nsew signal input
rlabel metal2 s 47030 119200 47086 120000 6 ALU_Sel1[1]
port 34 nsew signal input
rlabel metal2 s 29918 119200 29974 120000 6 ALU_Sel2[0]
port 35 nsew signal input
rlabel metal2 s 55678 119200 55734 120000 6 ALU_Sel2[1]
port 36 nsew signal input
rlabel metal3 s 179200 21360 180000 21480 6 B0[0]
port 37 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 B0[1]
port 38 nsew signal input
rlabel metal3 s 179200 64200 180000 64320 6 B0[2]
port 39 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 B0[3]
port 40 nsew signal input
rlabel metal2 s 107106 119200 107162 120000 6 B0[4]
port 41 nsew signal input
rlabel metal3 s 179200 98472 180000 98592 6 B0[5]
port 42 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 B0[6]
port 43 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 B0[7]
port 44 nsew signal input
rlabel metal3 s 179200 29928 180000 30048 6 B1[0]
port 45 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 B1[1]
port 46 nsew signal input
rlabel metal2 s 81346 119200 81402 120000 6 B1[2]
port 47 nsew signal input
rlabel metal2 s 89902 119200 89958 120000 6 B1[3]
port 48 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 B1[4]
port 49 nsew signal input
rlabel metal2 s 132774 119200 132830 120000 6 B1[5]
port 50 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 B1[6]
port 51 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 B1[7]
port 52 nsew signal input
rlabel metal2 s 4250 119200 4306 120000 6 CarryOut1
port 53 nsew signal output
rlabel metal3 s 179200 4224 180000 4344 6 CarryOut2
port 54 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 clk
port 55 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 57 nsew ground input
rlabel metal2 s 38474 119200 38530 120000 6 x[0]
port 58 nsew signal output
rlabel metal3 s 179200 47064 180000 47184 6 x[1]
port 59 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 x[2]
port 60 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 x[3]
port 61 nsew signal output
rlabel metal3 s 179200 89904 180000 90024 6 x[4]
port 62 nsew signal output
rlabel metal2 s 141422 119200 141478 120000 6 x[5]
port 63 nsew signal output
rlabel metal3 s 0 103504 800 103624 6 x[6]
port 64 nsew signal output
rlabel metal3 s 0 114384 800 114504 6 x[7]
port 65 nsew signal output
rlabel metal2 s 12806 119200 12862 120000 6 y
port 66 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6595250
string GDS_FILE /opt/caravel/caravel_example/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 421852
<< end >>

