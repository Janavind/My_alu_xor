magic
tech sky130A
magscale 1 2
timestamp 1647273520
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 1844 178848 117552
<< metal2 >>
rect 7470 119200 7526 120000
rect 22466 119200 22522 120000
rect 37462 119200 37518 120000
rect 52458 119200 52514 120000
rect 67454 119200 67510 120000
rect 82450 119200 82506 120000
rect 97446 119200 97502 120000
rect 112442 119200 112498 120000
rect 127438 119200 127494 120000
rect 142434 119200 142490 120000
rect 157430 119200 157486 120000
rect 172426 119200 172482 120000
rect 4986 0 5042 800
rect 14922 0 14978 800
rect 24950 0 25006 800
rect 34978 0 35034 800
rect 44914 0 44970 800
rect 54942 0 54998 800
rect 64970 0 65026 800
rect 74998 0 75054 800
rect 84934 0 84990 800
rect 94962 0 95018 800
rect 104990 0 105046 800
rect 114926 0 114982 800
rect 124954 0 125010 800
rect 134982 0 135038 800
rect 145010 0 145066 800
rect 154946 0 155002 800
rect 164974 0 165030 800
rect 175002 0 175058 800
<< obsm2 >>
rect 1398 119144 7414 119354
rect 7582 119144 22410 119354
rect 22578 119144 37406 119354
rect 37574 119144 52402 119354
rect 52570 119144 67398 119354
rect 67566 119144 82394 119354
rect 82562 119144 97390 119354
rect 97558 119144 112386 119354
rect 112554 119144 127382 119354
rect 127550 119144 142378 119354
rect 142546 119144 157374 119354
rect 157542 119144 172370 119354
rect 172538 119144 178186 119354
rect 1398 856 178186 119144
rect 1398 800 4930 856
rect 5098 800 14866 856
rect 15034 800 24894 856
rect 25062 800 34922 856
rect 35090 800 44858 856
rect 45026 800 54886 856
rect 55054 800 64914 856
rect 65082 800 74942 856
rect 75110 800 84878 856
rect 85046 800 94906 856
rect 95074 800 104934 856
rect 105102 800 114870 856
rect 115038 800 124898 856
rect 125066 800 134926 856
rect 135094 800 144954 856
rect 145122 800 154890 856
rect 155058 800 164918 856
rect 165086 800 174946 856
rect 175114 800 178186 856
<< metal3 >>
rect 179200 116696 180000 116816
rect 0 115880 800 116000
rect 179200 110440 180000 110560
rect 0 107856 800 107976
rect 179200 104048 180000 104168
rect 0 99832 800 99952
rect 179200 97792 180000 97912
rect 0 91808 800 91928
rect 179200 91400 180000 91520
rect 179200 85144 180000 85264
rect 0 83920 800 84040
rect 179200 78888 180000 79008
rect 0 75896 800 76016
rect 179200 72496 180000 72616
rect 0 67872 800 67992
rect 179200 66240 180000 66360
rect 0 59848 800 59968
rect 179200 59848 180000 59968
rect 179200 53592 180000 53712
rect 0 51824 800 51944
rect 179200 47200 180000 47320
rect 0 43936 800 44056
rect 179200 40944 180000 41064
rect 0 35912 800 36032
rect 179200 34688 180000 34808
rect 179200 28296 180000 28416
rect 0 27888 800 28008
rect 179200 22040 180000 22160
rect 0 19864 800 19984
rect 179200 15648 180000 15768
rect 0 11840 800 11960
rect 179200 9392 180000 9512
rect 0 3952 800 4072
rect 179200 3136 180000 3256
<< obsm3 >>
rect 800 116896 179200 117537
rect 800 116616 179120 116896
rect 800 116080 179200 116616
rect 880 115800 179200 116080
rect 800 110640 179200 115800
rect 800 110360 179120 110640
rect 800 108056 179200 110360
rect 880 107776 179200 108056
rect 800 104248 179200 107776
rect 800 103968 179120 104248
rect 800 100032 179200 103968
rect 880 99752 179200 100032
rect 800 97992 179200 99752
rect 800 97712 179120 97992
rect 800 92008 179200 97712
rect 880 91728 179200 92008
rect 800 91600 179200 91728
rect 800 91320 179120 91600
rect 800 85344 179200 91320
rect 800 85064 179120 85344
rect 800 84120 179200 85064
rect 880 83840 179200 84120
rect 800 79088 179200 83840
rect 800 78808 179120 79088
rect 800 76096 179200 78808
rect 880 75816 179200 76096
rect 800 72696 179200 75816
rect 800 72416 179120 72696
rect 800 68072 179200 72416
rect 880 67792 179200 68072
rect 800 66440 179200 67792
rect 800 66160 179120 66440
rect 800 60048 179200 66160
rect 880 59768 179120 60048
rect 800 53792 179200 59768
rect 800 53512 179120 53792
rect 800 52024 179200 53512
rect 880 51744 179200 52024
rect 800 47400 179200 51744
rect 800 47120 179120 47400
rect 800 44136 179200 47120
rect 880 43856 179200 44136
rect 800 41144 179200 43856
rect 800 40864 179120 41144
rect 800 36112 179200 40864
rect 880 35832 179200 36112
rect 800 34888 179200 35832
rect 800 34608 179120 34888
rect 800 28496 179200 34608
rect 800 28216 179120 28496
rect 800 28088 179200 28216
rect 880 27808 179200 28088
rect 800 22240 179200 27808
rect 800 21960 179120 22240
rect 800 20064 179200 21960
rect 880 19784 179200 20064
rect 800 15848 179200 19784
rect 800 15568 179120 15848
rect 800 12040 179200 15568
rect 880 11760 179200 12040
rect 800 9592 179200 11760
rect 800 9312 179120 9592
rect 800 4152 179200 9312
rect 880 3872 179200 4152
rect 800 3336 179200 3872
rect 800 3056 179120 3336
rect 800 2143 179200 3056
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 92979 3435 96288 65109
rect 96768 3435 100589 65109
<< labels >>
rlabel metal2 s 14922 0 14978 800 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 A0[2]
port 3 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 179200 85144 180000 85264 6 A0[5]
port 6 nsew signal input
rlabel metal2 s 112442 119200 112498 120000 6 A0[6]
port 7 nsew signal input
rlabel metal2 s 142434 119200 142490 120000 6 A0[7]
port 8 nsew signal input
rlabel metal2 s 7470 119200 7526 120000 6 A1[0]
port 9 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 A1[1]
port 10 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 A1[2]
port 11 nsew signal input
rlabel metal3 s 179200 66240 180000 66360 6 A1[3]
port 12 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 A1[4]
port 13 nsew signal input
rlabel metal2 s 67454 119200 67510 120000 6 A1[5]
port 14 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 A1[6]
port 15 nsew signal input
rlabel metal3 s 179200 116696 180000 116816 6 A1[7]
port 16 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 ALU_Out1[0]
port 17 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 ALU_Out1[1]
port 18 nsew signal output
rlabel metal3 s 0 51824 800 51944 6 ALU_Out1[2]
port 19 nsew signal output
rlabel metal3 s 179200 72496 180000 72616 6 ALU_Out1[3]
port 20 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 ALU_Out1[4]
port 21 nsew signal output
rlabel metal3 s 179200 91400 180000 91520 6 ALU_Out1[5]
port 22 nsew signal output
rlabel metal2 s 164974 0 165030 800 6 ALU_Out1[6]
port 23 nsew signal output
rlabel metal2 s 157430 119200 157486 120000 6 ALU_Out1[7]
port 24 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 ALU_Out2[0]
port 25 nsew signal output
rlabel metal2 s 22466 119200 22522 120000 6 ALU_Out2[1]
port 26 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 ALU_Out2[2]
port 27 nsew signal output
rlabel metal3 s 0 67872 800 67992 6 ALU_Out2[3]
port 28 nsew signal output
rlabel metal2 s 52458 119200 52514 120000 6 ALU_Out2[4]
port 29 nsew signal output
rlabel metal2 s 82450 119200 82506 120000 6 ALU_Out2[5]
port 30 nsew signal output
rlabel metal3 s 179200 104048 180000 104168 6 ALU_Out2[6]
port 31 nsew signal output
rlabel metal3 s 0 107856 800 107976 6 ALU_Out2[7]
port 32 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 ALU_Sel1[0]
port 33 nsew signal input
rlabel metal3 s 179200 34688 180000 34808 6 ALU_Sel1[1]
port 34 nsew signal input
rlabel metal3 s 179200 15648 180000 15768 6 ALU_Sel2[0]
port 35 nsew signal input
rlabel metal3 s 179200 40944 180000 41064 6 ALU_Sel2[1]
port 36 nsew signal input
rlabel metal3 s 179200 22040 180000 22160 6 B0[0]
port 37 nsew signal input
rlabel metal3 s 179200 47200 180000 47320 6 B0[1]
port 38 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 B0[2]
port 39 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 B0[3]
port 40 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 B0[4]
port 41 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 B0[5]
port 42 nsew signal input
rlabel metal3 s 179200 110440 180000 110560 6 B0[6]
port 43 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 B0[7]
port 44 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 B1[0]
port 45 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 B1[1]
port 46 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 B1[2]
port 47 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 B1[3]
port 48 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 B1[4]
port 49 nsew signal input
rlabel metal3 s 179200 97792 180000 97912 6 B1[5]
port 50 nsew signal input
rlabel metal2 s 127438 119200 127494 120000 6 B1[6]
port 51 nsew signal input
rlabel metal3 s 0 115880 800 116000 6 B1[7]
port 52 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 CarryOut1
port 53 nsew signal output
rlabel metal3 s 179200 3136 180000 3256 6 CarryOut2
port 54 nsew signal output
rlabel metal3 s 179200 9392 180000 9512 6 clk
port 55 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 57 nsew ground input
rlabel metal3 s 179200 28296 180000 28416 6 x[0]
port 58 nsew signal output
rlabel metal3 s 179200 53592 180000 53712 6 x[1]
port 59 nsew signal output
rlabel metal3 s 179200 59848 180000 59968 6 x[2]
port 60 nsew signal output
rlabel metal2 s 37462 119200 37518 120000 6 x[3]
port 61 nsew signal output
rlabel metal3 s 179200 78888 180000 79008 6 x[4]
port 62 nsew signal output
rlabel metal2 s 97446 119200 97502 120000 6 x[5]
port 63 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 x[6]
port 64 nsew signal output
rlabel metal2 s 172426 119200 172482 120000 6 x[7]
port 65 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 y
port 66 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6581092
string GDS_FILE /opt/caravel/caravel_example/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 417052
<< end >>

