magic
tech sky130A
magscale 1 2
timestamp 1647300040
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 7470 119200 7526 120000
rect 22466 119200 22522 120000
rect 37462 119200 37518 120000
rect 52458 119200 52514 120000
rect 67454 119200 67510 120000
rect 82450 119200 82506 120000
rect 97446 119200 97502 120000
rect 112442 119200 112498 120000
rect 127438 119200 127494 120000
rect 142434 119200 142490 120000
rect 157430 119200 157486 120000
rect 172426 119200 172482 120000
rect 5630 0 5686 800
rect 16854 0 16910 800
rect 28078 0 28134 800
rect 39302 0 39358 800
rect 50618 0 50674 800
rect 61842 0 61898 800
rect 73066 0 73122 800
rect 84382 0 84438 800
rect 95606 0 95662 800
rect 106830 0 106886 800
rect 118146 0 118202 800
rect 129370 0 129426 800
rect 140594 0 140650 800
rect 151910 0 151966 800
rect 163134 0 163190 800
rect 174358 0 174414 800
<< obsm2 >>
rect 1398 119144 7414 119354
rect 7582 119144 22410 119354
rect 22578 119144 37406 119354
rect 37574 119144 52402 119354
rect 52570 119144 67398 119354
rect 67566 119144 82394 119354
rect 82562 119144 97390 119354
rect 97558 119144 112386 119354
rect 112554 119144 127382 119354
rect 127550 119144 142378 119354
rect 142546 119144 157374 119354
rect 157542 119144 172370 119354
rect 172538 119144 178186 119354
rect 1398 856 178186 119144
rect 1398 800 5574 856
rect 5742 800 16798 856
rect 16966 800 28022 856
rect 28190 800 39246 856
rect 39414 800 50562 856
rect 50730 800 61786 856
rect 61954 800 73010 856
rect 73178 800 84326 856
rect 84494 800 95550 856
rect 95718 800 106774 856
rect 106942 800 118090 856
rect 118258 800 129314 856
rect 129482 800 140538 856
rect 140706 800 151854 856
rect 152022 800 163078 856
rect 163246 800 174302 856
rect 174470 800 178186 856
<< metal3 >>
rect 0 117104 800 117224
rect 179200 115880 180000 116000
rect 0 111392 800 111512
rect 179200 107856 180000 107976
rect 0 105680 800 105800
rect 0 99968 800 100088
rect 179200 99832 180000 99952
rect 0 94256 800 94376
rect 179200 91808 180000 91928
rect 0 88544 800 88664
rect 179200 83920 180000 84040
rect 0 82832 800 82952
rect 0 77120 800 77240
rect 179200 75896 180000 76016
rect 0 71408 800 71528
rect 179200 67872 180000 67992
rect 0 65696 800 65816
rect 0 59984 800 60104
rect 179200 59848 180000 59968
rect 0 54272 800 54392
rect 179200 51824 180000 51944
rect 0 48560 800 48680
rect 179200 43936 180000 44056
rect 0 42848 800 42968
rect 0 37136 800 37256
rect 179200 35912 180000 36032
rect 0 31424 800 31544
rect 179200 27888 180000 28008
rect 0 25712 800 25832
rect 0 20000 800 20120
rect 179200 19864 180000 19984
rect 0 14288 800 14408
rect 179200 11840 180000 11960
rect 0 8576 800 8696
rect 179200 3952 180000 4072
rect 0 2864 800 2984
<< obsm3 >>
rect 800 117304 179200 117537
rect 880 117024 179200 117304
rect 800 116080 179200 117024
rect 800 115800 179120 116080
rect 800 111592 179200 115800
rect 880 111312 179200 111592
rect 800 108056 179200 111312
rect 800 107776 179120 108056
rect 800 105880 179200 107776
rect 880 105600 179200 105880
rect 800 100168 179200 105600
rect 880 100032 179200 100168
rect 880 99888 179120 100032
rect 800 99752 179120 99888
rect 800 94456 179200 99752
rect 880 94176 179200 94456
rect 800 92008 179200 94176
rect 800 91728 179120 92008
rect 800 88744 179200 91728
rect 880 88464 179200 88744
rect 800 84120 179200 88464
rect 800 83840 179120 84120
rect 800 83032 179200 83840
rect 880 82752 179200 83032
rect 800 77320 179200 82752
rect 880 77040 179200 77320
rect 800 76096 179200 77040
rect 800 75816 179120 76096
rect 800 71608 179200 75816
rect 880 71328 179200 71608
rect 800 68072 179200 71328
rect 800 67792 179120 68072
rect 800 65896 179200 67792
rect 880 65616 179200 65896
rect 800 60184 179200 65616
rect 880 60048 179200 60184
rect 880 59904 179120 60048
rect 800 59768 179120 59904
rect 800 54472 179200 59768
rect 880 54192 179200 54472
rect 800 52024 179200 54192
rect 800 51744 179120 52024
rect 800 48760 179200 51744
rect 880 48480 179200 48760
rect 800 44136 179200 48480
rect 800 43856 179120 44136
rect 800 43048 179200 43856
rect 880 42768 179200 43048
rect 800 37336 179200 42768
rect 880 37056 179200 37336
rect 800 36112 179200 37056
rect 800 35832 179120 36112
rect 800 31624 179200 35832
rect 880 31344 179200 31624
rect 800 28088 179200 31344
rect 800 27808 179120 28088
rect 800 25912 179200 27808
rect 880 25632 179200 25912
rect 800 20200 179200 25632
rect 880 20064 179200 20200
rect 880 19920 179120 20064
rect 800 19784 179120 19920
rect 800 14488 179200 19784
rect 880 14208 179200 14488
rect 800 12040 179200 14208
rect 800 11760 179120 12040
rect 800 8776 179200 11760
rect 880 8496 179200 8776
rect 800 4152 179200 8496
rect 800 3872 179120 4152
rect 800 3064 179200 3872
rect 880 2784 179200 3064
rect 800 2143 179200 2784
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 75867 20435 80928 62797
rect 81408 20435 83661 62797
<< labels >>
rlabel metal2 s 22466 119200 22522 120000 6 A0[0]
port 1 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 0 31424 800 31544 6 A0[2]
port 3 nsew signal input
rlabel metal2 s 52458 119200 52514 120000 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 0 94256 800 94376 6 A0[5]
port 6 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 A0[6]
port 7 nsew signal input
rlabel metal2 s 127438 119200 127494 120000 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 A1[0]
port 9 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 A1[1]
port 10 nsew signal input
rlabel metal3 s 179200 51824 180000 51944 6 A1[2]
port 11 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 A1[3]
port 12 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 A1[4]
port 13 nsew signal input
rlabel metal2 s 97446 119200 97502 120000 6 A1[5]
port 14 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 A1[6]
port 15 nsew signal input
rlabel metal3 s 179200 107856 180000 107976 6 A1[7]
port 16 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 ALU_Out1[0]
port 17 nsew signal output
rlabel metal3 s 179200 27888 180000 28008 6 ALU_Out1[1]
port 18 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 ALU_Out1[2]
port 19 nsew signal output
rlabel metal3 s 179200 67872 180000 67992 6 ALU_Out1[3]
port 20 nsew signal output
rlabel metal3 s 0 77120 800 77240 6 ALU_Out1[4]
port 21 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 ALU_Out1[5]
port 22 nsew signal output
rlabel metal2 s 140594 0 140650 800 6 ALU_Out1[6]
port 23 nsew signal output
rlabel metal3 s 179200 115880 180000 116000 6 ALU_Out1[7]
port 24 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 ALU_Out2[0]
port 25 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 ALU_Out2[1]
port 26 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 ALU_Out2[2]
port 27 nsew signal output
rlabel metal3 s 179200 75896 180000 76016 6 ALU_Out2[3]
port 28 nsew signal output
rlabel metal3 s 179200 83920 180000 84040 6 ALU_Out2[4]
port 29 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 ALU_Out2[5]
port 30 nsew signal output
rlabel metal2 s 112442 119200 112498 120000 6 ALU_Out2[6]
port 31 nsew signal output
rlabel metal2 s 142434 119200 142490 120000 6 ALU_Out2[7]
port 32 nsew signal output
rlabel metal3 s 179200 11840 180000 11960 6 ALU_Sel1[0]
port 33 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 ALU_Sel1[1]
port 34 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 ALU_Sel2[0]
port 35 nsew signal input
rlabel metal3 s 179200 35912 180000 36032 6 ALU_Sel2[1]
port 36 nsew signal input
rlabel metal3 s 179200 19864 180000 19984 6 B0[0]
port 37 nsew signal input
rlabel metal3 s 179200 43936 180000 44056 6 B0[1]
port 38 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 B0[2]
port 39 nsew signal input
rlabel metal2 s 67454 119200 67510 120000 6 B0[3]
port 40 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 B0[4]
port 41 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 B0[5]
port 42 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 B0[6]
port 43 nsew signal input
rlabel metal2 s 157430 119200 157486 120000 6 B0[7]
port 44 nsew signal input
rlabel metal2 s 37462 119200 37518 120000 6 B1[0]
port 45 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 B1[1]
port 46 nsew signal input
rlabel metal3 s 179200 59848 180000 59968 6 B1[2]
port 47 nsew signal input
rlabel metal2 s 82450 119200 82506 120000 6 B1[3]
port 48 nsew signal input
rlabel metal3 s 179200 91808 180000 91928 6 B1[4]
port 49 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 B1[5]
port 50 nsew signal input
rlabel metal3 s 179200 99832 180000 99952 6 B1[6]
port 51 nsew signal input
rlabel metal2 s 172426 119200 172482 120000 6 B1[7]
port 52 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 CarryOut1
port 53 nsew signal output
rlabel metal2 s 7470 119200 7526 120000 6 CarryOut2
port 54 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 clk
port 55 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 57 nsew ground input
rlabel metal2 s 39302 0 39358 800 6 x[0]
port 58 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 x[1]
port 59 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 x[2]
port 60 nsew signal output
rlabel metal3 s 0 59984 800 60104 6 x[3]
port 61 nsew signal output
rlabel metal3 s 0 88544 800 88664 6 x[4]
port 62 nsew signal output
rlabel metal3 s 0 111392 800 111512 6 x[5]
port 63 nsew signal output
rlabel metal2 s 163134 0 163190 800 6 x[6]
port 64 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 x[7]
port 65 nsew signal output
rlabel metal3 s 179200 3952 180000 4072 6 y
port 66 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6559612
string GDS_FILE /opt/caravel/caravel_example/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 383476
<< end >>

