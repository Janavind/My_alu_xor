VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 404.640 900.000 405.240 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 596.000 750.170 600.000 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.720 4.000 511.320 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 17.040 900.000 17.640 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 157.800 900.000 158.400 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 546.080 900.000 546.680 ;
    END
  END A1[7]
  PIN ALU_Out1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END ALU_Out1[0]
  PIN ALU_Out1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END ALU_Out1[1]
  PIN ALU_Out1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 596.000 330.190 600.000 ;
    END
  END ALU_Out1[2]
  PIN ALU_Out1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END ALU_Out1[3]
  PIN ALU_Out1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 333.920 900.000 334.520 ;
    END
  END ALU_Out1[4]
  PIN ALU_Out1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 596.000 630.110 600.000 ;
    END
  END ALU_Out1[5]
  PIN ALU_Out1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 475.360 900.000 475.960 ;
    END
  END ALU_Out1[6]
  PIN ALU_Out1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 596.000 870.230 600.000 ;
    END
  END ALU_Out1[7]
  PIN ALU_Out2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 596.000 149.870 600.000 ;
    END
  END ALU_Out2[0]
  PIN ALU_Out2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END ALU_Out2[1]
  PIN ALU_Out2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 596.000 389.990 600.000 ;
    END
  END ALU_Out2[2]
  PIN ALU_Out2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 228.520 900.000 229.120 ;
    END
  END ALU_Out2[3]
  PIN ALU_Out2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END ALU_Out2[4]
  PIN ALU_Out2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 596.000 690.370 600.000 ;
    END
  END ALU_Out2[5]
  PIN ALU_Out2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 596.000 810.430 600.000 ;
    END
  END ALU_Out2[6]
  PIN ALU_Out2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 581.440 900.000 582.040 ;
    END
  END ALU_Out2[7]
  PIN ALU_Sel1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END ALU_Sel1[0]
  PIN ALU_Sel1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 122.440 900.000 123.040 ;
    END
  END ALU_Sel1[1]
  PIN ALU_Sel2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 51.720 900.000 52.320 ;
    END
  END ALU_Sel2[0]
  PIN ALU_Sel2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END ALU_Sel2[1]
  PIN B0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 87.080 900.000 87.680 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 596.000 269.930 600.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 596.000 450.250 600.000 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 263.880 900.000 264.480 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 369.280 900.000 369.880 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 596.000 210.130 600.000 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 596.000 510.050 600.000 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 299.240 900.000 299.840 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 475.360 4.000 475.960 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 0.000 870.230 4.000 ;
    END
  END B1[7]
  PIN CarryOut1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 596.000 30.270 600.000 ;
    END
  END CarryOut1
  PIN CarryOut2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 596.000 90.070 600.000 ;
    END
  END CarryOut2
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END clk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 193.160 900.000 193.760 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 596.000 570.310 600.000 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 440.000 900.000 440.600 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 510.720 900.000 511.320 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END x[7]
  PIN y
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END y
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 6.990 595.720 29.710 596.770 ;
        RECT 30.550 595.720 89.510 596.770 ;
        RECT 90.350 595.720 149.310 596.770 ;
        RECT 150.150 595.720 209.570 596.770 ;
        RECT 210.410 595.720 269.370 596.770 ;
        RECT 270.210 595.720 329.630 596.770 ;
        RECT 330.470 595.720 389.430 596.770 ;
        RECT 390.270 595.720 449.690 596.770 ;
        RECT 450.530 595.720 509.490 596.770 ;
        RECT 510.330 595.720 569.750 596.770 ;
        RECT 570.590 595.720 629.550 596.770 ;
        RECT 630.390 595.720 689.810 596.770 ;
        RECT 690.650 595.720 749.610 596.770 ;
        RECT 750.450 595.720 809.870 596.770 ;
        RECT 810.710 595.720 869.670 596.770 ;
        RECT 870.510 595.720 890.930 596.770 ;
        RECT 6.990 4.280 890.930 595.720 ;
        RECT 6.990 4.000 29.710 4.280 ;
        RECT 30.550 4.000 89.510 4.280 ;
        RECT 90.350 4.000 149.310 4.280 ;
        RECT 150.150 4.000 209.570 4.280 ;
        RECT 210.410 4.000 269.370 4.280 ;
        RECT 270.210 4.000 329.630 4.280 ;
        RECT 330.470 4.000 389.430 4.280 ;
        RECT 390.270 4.000 449.690 4.280 ;
        RECT 450.530 4.000 509.490 4.280 ;
        RECT 510.330 4.000 569.750 4.280 ;
        RECT 570.590 4.000 629.550 4.280 ;
        RECT 630.390 4.000 689.810 4.280 ;
        RECT 690.650 4.000 749.610 4.280 ;
        RECT 750.450 4.000 809.870 4.280 ;
        RECT 810.710 4.000 869.670 4.280 ;
        RECT 870.510 4.000 890.930 4.280 ;
      LAYER met3 ;
        RECT 4.000 582.440 896.000 587.685 ;
        RECT 4.400 581.040 895.600 582.440 ;
        RECT 4.000 547.080 896.000 581.040 ;
        RECT 4.400 545.680 895.600 547.080 ;
        RECT 4.000 511.720 896.000 545.680 ;
        RECT 4.400 510.320 895.600 511.720 ;
        RECT 4.000 476.360 896.000 510.320 ;
        RECT 4.400 474.960 895.600 476.360 ;
        RECT 4.000 441.000 896.000 474.960 ;
        RECT 4.400 439.600 895.600 441.000 ;
        RECT 4.000 405.640 896.000 439.600 ;
        RECT 4.400 404.240 895.600 405.640 ;
        RECT 4.000 370.280 896.000 404.240 ;
        RECT 4.400 368.880 895.600 370.280 ;
        RECT 4.000 334.920 896.000 368.880 ;
        RECT 4.400 333.520 895.600 334.920 ;
        RECT 4.000 300.240 896.000 333.520 ;
        RECT 4.400 298.840 895.600 300.240 ;
        RECT 4.000 264.880 896.000 298.840 ;
        RECT 4.400 263.480 895.600 264.880 ;
        RECT 4.000 229.520 896.000 263.480 ;
        RECT 4.400 228.120 895.600 229.520 ;
        RECT 4.000 194.160 896.000 228.120 ;
        RECT 4.400 192.760 895.600 194.160 ;
        RECT 4.000 158.800 896.000 192.760 ;
        RECT 4.400 157.400 895.600 158.800 ;
        RECT 4.000 123.440 896.000 157.400 ;
        RECT 4.400 122.040 895.600 123.440 ;
        RECT 4.000 88.080 896.000 122.040 ;
        RECT 4.400 86.680 895.600 88.080 ;
        RECT 4.000 52.720 896.000 86.680 ;
        RECT 4.400 51.320 895.600 52.720 ;
        RECT 4.000 18.040 896.000 51.320 ;
        RECT 4.400 16.640 895.600 18.040 ;
        RECT 4.000 10.715 896.000 16.640 ;
      LAYER met4 ;
        RECT 437.295 273.535 480.865 373.825 ;
  END
END user_proj_example
END LIBRARY

