magic
tech sky130A
magscale 1 2
timestamp 1647279819
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 5998 119200 6054 120000
rect 17958 119200 18014 120000
rect 29918 119200 29974 120000
rect 41970 119200 42026 120000
rect 53930 119200 53986 120000
rect 65982 119200 66038 120000
rect 77942 119200 77998 120000
rect 89994 119200 90050 120000
rect 101954 119200 102010 120000
rect 114006 119200 114062 120000
rect 125966 119200 126022 120000
rect 138018 119200 138074 120000
rect 149978 119200 150034 120000
rect 162030 119200 162086 120000
rect 173990 119200 174046 120000
rect 5998 0 6054 800
rect 17958 0 18014 800
rect 29918 0 29974 800
rect 41970 0 42026 800
rect 53930 0 53986 800
rect 65982 0 66038 800
rect 77942 0 77998 800
rect 89994 0 90050 800
rect 101954 0 102010 800
rect 114006 0 114062 800
rect 125966 0 126022 800
rect 138018 0 138074 800
rect 149978 0 150034 800
rect 162030 0 162086 800
rect 173990 0 174046 800
<< obsm2 >>
rect 1398 119144 5942 119354
rect 6110 119144 17902 119354
rect 18070 119144 29862 119354
rect 30030 119144 41914 119354
rect 42082 119144 53874 119354
rect 54042 119144 65926 119354
rect 66094 119144 77886 119354
rect 78054 119144 89938 119354
rect 90106 119144 101898 119354
rect 102066 119144 113950 119354
rect 114118 119144 125910 119354
rect 126078 119144 137962 119354
rect 138130 119144 149922 119354
rect 150090 119144 161974 119354
rect 162142 119144 173934 119354
rect 174102 119144 178186 119354
rect 1398 856 178186 119144
rect 1398 800 5942 856
rect 6110 800 17902 856
rect 18070 800 29862 856
rect 30030 800 41914 856
rect 42082 800 53874 856
rect 54042 800 65926 856
rect 66094 800 77886 856
rect 78054 800 89938 856
rect 90106 800 101898 856
rect 102066 800 113950 856
rect 114118 800 125910 856
rect 126078 800 137962 856
rect 138130 800 149922 856
rect 150090 800 161974 856
rect 162142 800 173934 856
rect 174102 800 178186 856
<< metal3 >>
rect 0 116288 800 116408
rect 179200 116288 180000 116408
rect 0 109216 800 109336
rect 179200 109216 180000 109336
rect 0 102144 800 102264
rect 179200 102144 180000 102264
rect 0 95072 800 95192
rect 179200 95072 180000 95192
rect 0 88000 800 88120
rect 179200 88000 180000 88120
rect 0 80928 800 81048
rect 179200 80928 180000 81048
rect 0 73856 800 73976
rect 179200 73856 180000 73976
rect 0 66784 800 66904
rect 179200 66784 180000 66904
rect 0 59848 800 59968
rect 179200 59848 180000 59968
rect 0 52776 800 52896
rect 179200 52776 180000 52896
rect 0 45704 800 45824
rect 179200 45704 180000 45824
rect 0 38632 800 38752
rect 179200 38632 180000 38752
rect 0 31560 800 31680
rect 179200 31560 180000 31680
rect 0 24488 800 24608
rect 179200 24488 180000 24608
rect 0 17416 800 17536
rect 179200 17416 180000 17536
rect 0 10344 800 10464
rect 179200 10344 180000 10464
rect 0 3408 800 3528
rect 179200 3408 180000 3528
<< obsm3 >>
rect 800 116488 179200 117537
rect 880 116208 179120 116488
rect 800 109416 179200 116208
rect 880 109136 179120 109416
rect 800 102344 179200 109136
rect 880 102064 179120 102344
rect 800 95272 179200 102064
rect 880 94992 179120 95272
rect 800 88200 179200 94992
rect 880 87920 179120 88200
rect 800 81128 179200 87920
rect 880 80848 179120 81128
rect 800 74056 179200 80848
rect 880 73776 179120 74056
rect 800 66984 179200 73776
rect 880 66704 179120 66984
rect 800 60048 179200 66704
rect 880 59768 179120 60048
rect 800 52976 179200 59768
rect 880 52696 179120 52976
rect 800 45904 179200 52696
rect 880 45624 179120 45904
rect 800 38832 179200 45624
rect 880 38552 179120 38832
rect 800 31760 179200 38552
rect 880 31480 179120 31760
rect 800 24688 179200 31480
rect 880 24408 179120 24688
rect 800 17616 179200 24408
rect 880 17336 179120 17616
rect 800 10544 179200 17336
rect 880 10264 179120 10544
rect 800 3608 179200 10264
rect 880 3328 179120 3608
rect 800 2143 179200 3328
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 87459 54707 96173 74765
<< labels >>
rlabel metal2 s 17958 0 18014 800 6 A0[0]
port 1 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 A0[1]
port 2 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 179200 80928 180000 81048 6 A0[5]
port 6 nsew signal input
rlabel metal2 s 149978 119200 150034 120000 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 0 102144 800 102264 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 179200 3408 180000 3528 6 A1[0]
port 9 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 A1[1]
port 10 nsew signal input
rlabel metal3 s 179200 31560 180000 31680 6 A1[2]
port 11 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 A1[3]
port 12 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 A1[4]
port 13 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 A1[5]
port 14 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 A1[6]
port 15 nsew signal input
rlabel metal3 s 179200 109216 180000 109336 6 A1[7]
port 16 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 ALU_Out1[0]
port 17 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 ALU_Out1[1]
port 18 nsew signal output
rlabel metal2 s 65982 119200 66038 120000 6 ALU_Out1[2]
port 19 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 ALU_Out1[3]
port 20 nsew signal output
rlabel metal3 s 179200 66784 180000 66904 6 ALU_Out1[4]
port 21 nsew signal output
rlabel metal2 s 125966 119200 126022 120000 6 ALU_Out1[5]
port 22 nsew signal output
rlabel metal3 s 179200 95072 180000 95192 6 ALU_Out1[6]
port 23 nsew signal output
rlabel metal2 s 173990 119200 174046 120000 6 ALU_Out1[7]
port 24 nsew signal output
rlabel metal2 s 29918 119200 29974 120000 6 ALU_Out2[0]
port 25 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 ALU_Out2[1]
port 26 nsew signal output
rlabel metal2 s 77942 119200 77998 120000 6 ALU_Out2[2]
port 27 nsew signal output
rlabel metal3 s 179200 45704 180000 45824 6 ALU_Out2[3]
port 28 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 ALU_Out2[4]
port 29 nsew signal output
rlabel metal2 s 138018 119200 138074 120000 6 ALU_Out2[5]
port 30 nsew signal output
rlabel metal2 s 162030 119200 162086 120000 6 ALU_Out2[6]
port 31 nsew signal output
rlabel metal3 s 179200 116288 180000 116408 6 ALU_Out2[7]
port 32 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 ALU_Sel1[0]
port 33 nsew signal input
rlabel metal3 s 179200 24488 180000 24608 6 ALU_Sel1[1]
port 34 nsew signal input
rlabel metal3 s 179200 10344 180000 10464 6 ALU_Sel2[0]
port 35 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 ALU_Sel2[1]
port 36 nsew signal input
rlabel metal3 s 179200 17416 180000 17536 6 B0[0]
port 37 nsew signal input
rlabel metal2 s 53930 119200 53986 120000 6 B0[1]
port 38 nsew signal input
rlabel metal2 s 89994 119200 90050 120000 6 B0[2]
port 39 nsew signal input
rlabel metal3 s 179200 52776 180000 52896 6 B0[3]
port 40 nsew signal input
rlabel metal3 s 179200 73856 180000 73976 6 B0[4]
port 41 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 B0[5]
port 42 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 B0[6]
port 43 nsew signal input
rlabel metal3 s 0 109216 800 109336 6 B0[7]
port 44 nsew signal input
rlabel metal2 s 41970 119200 42026 120000 6 B1[0]
port 45 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 B1[1]
port 46 nsew signal input
rlabel metal2 s 101954 119200 102010 120000 6 B1[2]
port 47 nsew signal input
rlabel metal3 s 179200 59848 180000 59968 6 B1[3]
port 48 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 B1[4]
port 49 nsew signal input
rlabel metal3 s 0 95072 800 95192 6 B1[5]
port 50 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 B1[6]
port 51 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 B1[7]
port 52 nsew signal input
rlabel metal2 s 5998 119200 6054 120000 6 CarryOut1
port 53 nsew signal output
rlabel metal2 s 17958 119200 18014 120000 6 CarryOut2
port 54 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 clk
port 55 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 57 nsew ground input
rlabel metal3 s 0 24488 800 24608 6 x[0]
port 58 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 x[1]
port 59 nsew signal output
rlabel metal3 s 179200 38632 180000 38752 6 x[2]
port 60 nsew signal output
rlabel metal2 s 114006 119200 114062 120000 6 x[3]
port 61 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 x[4]
port 62 nsew signal output
rlabel metal3 s 179200 88000 180000 88120 6 x[5]
port 63 nsew signal output
rlabel metal3 s 179200 102144 180000 102264 6 x[6]
port 64 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 x[7]
port 65 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 y
port 66 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6779538
string GDS_FILE /opt/caravel/caravel_example/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 495082
<< end >>

