VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 192.480 900.000 193.080 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 596.000 321.450 600.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 363.840 900.000 364.440 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 596.000 750.170 600.000 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 4.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 596.000 364.230 600.000 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 596.000 578.590 600.000 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 596.000 835.730 600.000 ;
    END
  END A1[7]
  PIN ALU_Out1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END ALU_Out1[0]
  PIN ALU_Out1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END ALU_Out1[1]
  PIN ALU_Out1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 278.160 900.000 278.760 ;
    END
  END ALU_Out1[2]
  PIN ALU_Out1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END ALU_Out1[3]
  PIN ALU_Out1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 596.000 493.030 600.000 ;
    END
  END ALU_Out1[4]
  PIN ALU_Out1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 596.000 621.370 600.000 ;
    END
  END ALU_Out1[5]
  PIN ALU_Out1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 596.000 792.950 600.000 ;
    END
  END ALU_Out1[6]
  PIN ALU_Out1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.230 596.000 878.510 600.000 ;
    END
  END ALU_Out1[7]
  PIN ALU_Out2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 596.000 107.090 600.000 ;
    END
  END ALU_Out2[0]
  PIN ALU_Out2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END ALU_Out2[1]
  PIN ALU_Out2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END ALU_Out2[2]
  PIN ALU_Out2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END ALU_Out2[3]
  PIN ALU_Out2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 406.680 900.000 407.280 ;
    END
  END ALU_Out2[4]
  PIN ALU_Out2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END ALU_Out2[5]
  PIN ALU_Out2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 535.200 900.000 535.800 ;
    END
  END ALU_Out2[6]
  PIN ALU_Out2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 578.040 900.000 578.640 ;
    END
  END ALU_Out2[7]
  PIN ALU_Sel1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 63.960 900.000 64.560 ;
    END
  END ALU_Sel1[0]
  PIN ALU_Sel1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 596.000 235.430 600.000 ;
    END
  END ALU_Sel1[1]
  PIN ALU_Sel2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 596.000 149.870 600.000 ;
    END
  END ALU_Sel2[0]
  PIN ALU_Sel2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 596.000 278.670 600.000 ;
    END
  END ALU_Sel2[1]
  PIN B0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 106.800 900.000 107.400 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 321.000 900.000 321.600 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 596.000 535.810 600.000 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 492.360 900.000 492.960 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 149.640 900.000 150.240 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 596.000 407.010 600.000 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 596.000 449.790 600.000 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 596.000 664.150 600.000 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END B1[7]
  PIN CarryOut1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 596.000 21.530 600.000 ;
    END
  END CarryOut1
  PIN CarryOut2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 21.120 900.000 21.720 ;
    END
  END CarryOut2
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END clk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 596.000 192.650 600.000 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 235.320 900.000 235.920 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 449.520 900.000 450.120 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 596.000 707.390 600.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END x[7]
  PIN y
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 596.000 64.310 600.000 ;
    END
  END y
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 9.560 894.240 587.760 ;
      LAYER met2 ;
        RECT 6.990 595.720 20.970 596.770 ;
        RECT 21.810 595.720 63.750 596.770 ;
        RECT 64.590 595.720 106.530 596.770 ;
        RECT 107.370 595.720 149.310 596.770 ;
        RECT 150.150 595.720 192.090 596.770 ;
        RECT 192.930 595.720 234.870 596.770 ;
        RECT 235.710 595.720 278.110 596.770 ;
        RECT 278.950 595.720 320.890 596.770 ;
        RECT 321.730 595.720 363.670 596.770 ;
        RECT 364.510 595.720 406.450 596.770 ;
        RECT 407.290 595.720 449.230 596.770 ;
        RECT 450.070 595.720 492.470 596.770 ;
        RECT 493.310 595.720 535.250 596.770 ;
        RECT 536.090 595.720 578.030 596.770 ;
        RECT 578.870 595.720 620.810 596.770 ;
        RECT 621.650 595.720 663.590 596.770 ;
        RECT 664.430 595.720 706.830 596.770 ;
        RECT 707.670 595.720 749.610 596.770 ;
        RECT 750.450 595.720 792.390 596.770 ;
        RECT 793.230 595.720 835.170 596.770 ;
        RECT 836.010 595.720 877.950 596.770 ;
        RECT 878.790 595.720 890.930 596.770 ;
        RECT 6.990 4.280 890.930 595.720 ;
        RECT 6.990 4.000 24.650 4.280 ;
        RECT 25.490 4.000 74.330 4.280 ;
        RECT 75.170 4.000 124.470 4.280 ;
        RECT 125.310 4.000 174.610 4.280 ;
        RECT 175.450 4.000 224.290 4.280 ;
        RECT 225.130 4.000 274.430 4.280 ;
        RECT 275.270 4.000 324.570 4.280 ;
        RECT 325.410 4.000 374.710 4.280 ;
        RECT 375.550 4.000 424.390 4.280 ;
        RECT 425.230 4.000 474.530 4.280 ;
        RECT 475.370 4.000 524.670 4.280 ;
        RECT 525.510 4.000 574.350 4.280 ;
        RECT 575.190 4.000 624.490 4.280 ;
        RECT 625.330 4.000 674.630 4.280 ;
        RECT 675.470 4.000 724.770 4.280 ;
        RECT 725.610 4.000 774.450 4.280 ;
        RECT 775.290 4.000 824.590 4.280 ;
        RECT 825.430 4.000 874.730 4.280 ;
        RECT 875.570 4.000 890.930 4.280 ;
      LAYER met3 ;
        RECT 4.000 579.040 896.000 587.685 ;
        RECT 4.000 577.640 895.600 579.040 ;
        RECT 4.000 572.920 896.000 577.640 ;
        RECT 4.400 571.520 896.000 572.920 ;
        RECT 4.000 536.200 896.000 571.520 ;
        RECT 4.000 534.800 895.600 536.200 ;
        RECT 4.000 518.520 896.000 534.800 ;
        RECT 4.400 517.120 896.000 518.520 ;
        RECT 4.000 493.360 896.000 517.120 ;
        RECT 4.000 491.960 895.600 493.360 ;
        RECT 4.000 464.120 896.000 491.960 ;
        RECT 4.400 462.720 896.000 464.120 ;
        RECT 4.000 450.520 896.000 462.720 ;
        RECT 4.000 449.120 895.600 450.520 ;
        RECT 4.000 409.720 896.000 449.120 ;
        RECT 4.400 408.320 896.000 409.720 ;
        RECT 4.000 407.680 896.000 408.320 ;
        RECT 4.000 406.280 895.600 407.680 ;
        RECT 4.000 364.840 896.000 406.280 ;
        RECT 4.000 363.440 895.600 364.840 ;
        RECT 4.000 355.320 896.000 363.440 ;
        RECT 4.400 353.920 896.000 355.320 ;
        RECT 4.000 322.000 896.000 353.920 ;
        RECT 4.000 320.600 895.600 322.000 ;
        RECT 4.000 300.240 896.000 320.600 ;
        RECT 4.400 298.840 896.000 300.240 ;
        RECT 4.000 279.160 896.000 298.840 ;
        RECT 4.000 277.760 895.600 279.160 ;
        RECT 4.000 245.840 896.000 277.760 ;
        RECT 4.400 244.440 896.000 245.840 ;
        RECT 4.000 236.320 896.000 244.440 ;
        RECT 4.000 234.920 895.600 236.320 ;
        RECT 4.000 193.480 896.000 234.920 ;
        RECT 4.000 192.080 895.600 193.480 ;
        RECT 4.000 191.440 896.000 192.080 ;
        RECT 4.400 190.040 896.000 191.440 ;
        RECT 4.000 150.640 896.000 190.040 ;
        RECT 4.000 149.240 895.600 150.640 ;
        RECT 4.000 137.040 896.000 149.240 ;
        RECT 4.400 135.640 896.000 137.040 ;
        RECT 4.000 107.800 896.000 135.640 ;
        RECT 4.000 106.400 895.600 107.800 ;
        RECT 4.000 82.640 896.000 106.400 ;
        RECT 4.400 81.240 896.000 82.640 ;
        RECT 4.000 64.960 896.000 81.240 ;
        RECT 4.000 63.560 895.600 64.960 ;
        RECT 4.000 28.240 896.000 63.560 ;
        RECT 4.400 26.840 896.000 28.240 ;
        RECT 4.000 22.120 896.000 26.840 ;
        RECT 4.000 20.720 895.600 22.120 ;
        RECT 4.000 10.715 896.000 20.720 ;
      LAYER met4 ;
        RECT 447.415 23.295 481.440 376.545 ;
        RECT 483.840 23.295 498.345 376.545 ;
  END
END user_proj_example
END LIBRARY

