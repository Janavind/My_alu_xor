VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 425.720 900.000 426.320 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 596.000 562.490 600.000 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 596.000 712.450 600.000 ;
    END
  END A0[7]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 596.000 37.630 600.000 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 331.200 900.000 331.800 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 596.000 337.550 600.000 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 4.000 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 583.480 900.000 584.080 ;
    END
  END A1[7]
  PIN ALU_Out1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END ALU_Out1[0]
  PIN ALU_Out1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END ALU_Out1[1]
  PIN ALU_Out1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END ALU_Out1[2]
  PIN ALU_Out1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 362.480 900.000 363.080 ;
    END
  END ALU_Out1[3]
  PIN ALU_Out1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END ALU_Out1[4]
  PIN ALU_Out1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 457.000 900.000 457.600 ;
    END
  END ALU_Out1[5]
  PIN ALU_Out1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END ALU_Out1[6]
  PIN ALU_Out1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 596.000 787.430 600.000 ;
    END
  END ALU_Out1[7]
  PIN ALU_Out2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END ALU_Out2[0]
  PIN ALU_Out2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 596.000 112.610 600.000 ;
    END
  END ALU_Out2[1]
  PIN ALU_Out2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END ALU_Out2[2]
  PIN ALU_Out2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END ALU_Out2[3]
  PIN ALU_Out2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 596.000 262.570 600.000 ;
    END
  END ALU_Out2[4]
  PIN ALU_Out2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 596.000 412.530 600.000 ;
    END
  END ALU_Out2[5]
  PIN ALU_Out2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 520.240 900.000 520.840 ;
    END
  END ALU_Out2[6]
  PIN ALU_Out2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.280 4.000 539.880 ;
    END
  END ALU_Out2[7]
  PIN ALU_Sel1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END ALU_Sel1[0]
  PIN ALU_Sel1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 173.440 900.000 174.040 ;
    END
  END ALU_Sel1[1]
  PIN ALU_Sel2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 78.240 900.000 78.840 ;
    END
  END ALU_Sel2[0]
  PIN ALU_Sel2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 204.720 900.000 205.320 ;
    END
  END ALU_Sel2[1]
  PIN B0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 110.200 900.000 110.800 ;
    END
  END B0[0]
  PIN B0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 236.000 900.000 236.600 ;
    END
  END B0[1]
  PIN B0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END B0[2]
  PIN B0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END B0[3]
  PIN B0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END B0[4]
  PIN B0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END B0[5]
  PIN B0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 552.200 900.000 552.800 ;
    END
  END B0[6]
  PIN B0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END B0[7]
  PIN B1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END B1[0]
  PIN B1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END B1[1]
  PIN B1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END B1[2]
  PIN B1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END B1[3]
  PIN B1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END B1[4]
  PIN B1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 488.960 900.000 489.560 ;
    END
  END B1[5]
  PIN B1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 596.000 637.470 600.000 ;
    END
  END B1[6]
  PIN B1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END B1[7]
  PIN CarryOut1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END CarryOut1
  PIN CarryOut2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 15.680 900.000 16.280 ;
    END
  END CarryOut2
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 46.960 900.000 47.560 ;
    END
  END clk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 141.480 900.000 142.080 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 267.960 900.000 268.560 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 299.240 900.000 299.840 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 596.000 187.590 600.000 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 394.440 900.000 395.040 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 596.000 487.510 600.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 596.000 862.410 600.000 ;
    END
  END x[7]
  PIN y
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END y
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 9.220 894.240 587.760 ;
      LAYER met2 ;
        RECT 6.990 595.720 37.070 596.770 ;
        RECT 37.910 595.720 112.050 596.770 ;
        RECT 112.890 595.720 187.030 596.770 ;
        RECT 187.870 595.720 262.010 596.770 ;
        RECT 262.850 595.720 336.990 596.770 ;
        RECT 337.830 595.720 411.970 596.770 ;
        RECT 412.810 595.720 486.950 596.770 ;
        RECT 487.790 595.720 561.930 596.770 ;
        RECT 562.770 595.720 636.910 596.770 ;
        RECT 637.750 595.720 711.890 596.770 ;
        RECT 712.730 595.720 786.870 596.770 ;
        RECT 787.710 595.720 861.850 596.770 ;
        RECT 862.690 595.720 890.930 596.770 ;
        RECT 6.990 4.280 890.930 595.720 ;
        RECT 6.990 4.000 24.650 4.280 ;
        RECT 25.490 4.000 74.330 4.280 ;
        RECT 75.170 4.000 124.470 4.280 ;
        RECT 125.310 4.000 174.610 4.280 ;
        RECT 175.450 4.000 224.290 4.280 ;
        RECT 225.130 4.000 274.430 4.280 ;
        RECT 275.270 4.000 324.570 4.280 ;
        RECT 325.410 4.000 374.710 4.280 ;
        RECT 375.550 4.000 424.390 4.280 ;
        RECT 425.230 4.000 474.530 4.280 ;
        RECT 475.370 4.000 524.670 4.280 ;
        RECT 525.510 4.000 574.350 4.280 ;
        RECT 575.190 4.000 624.490 4.280 ;
        RECT 625.330 4.000 674.630 4.280 ;
        RECT 675.470 4.000 724.770 4.280 ;
        RECT 725.610 4.000 774.450 4.280 ;
        RECT 775.290 4.000 824.590 4.280 ;
        RECT 825.430 4.000 874.730 4.280 ;
        RECT 875.570 4.000 890.930 4.280 ;
      LAYER met3 ;
        RECT 4.000 584.480 896.000 587.685 ;
        RECT 4.000 583.080 895.600 584.480 ;
        RECT 4.000 580.400 896.000 583.080 ;
        RECT 4.400 579.000 896.000 580.400 ;
        RECT 4.000 553.200 896.000 579.000 ;
        RECT 4.000 551.800 895.600 553.200 ;
        RECT 4.000 540.280 896.000 551.800 ;
        RECT 4.400 538.880 896.000 540.280 ;
        RECT 4.000 521.240 896.000 538.880 ;
        RECT 4.000 519.840 895.600 521.240 ;
        RECT 4.000 500.160 896.000 519.840 ;
        RECT 4.400 498.760 896.000 500.160 ;
        RECT 4.000 489.960 896.000 498.760 ;
        RECT 4.000 488.560 895.600 489.960 ;
        RECT 4.000 460.040 896.000 488.560 ;
        RECT 4.400 458.640 896.000 460.040 ;
        RECT 4.000 458.000 896.000 458.640 ;
        RECT 4.000 456.600 895.600 458.000 ;
        RECT 4.000 426.720 896.000 456.600 ;
        RECT 4.000 425.320 895.600 426.720 ;
        RECT 4.000 420.600 896.000 425.320 ;
        RECT 4.400 419.200 896.000 420.600 ;
        RECT 4.000 395.440 896.000 419.200 ;
        RECT 4.000 394.040 895.600 395.440 ;
        RECT 4.000 380.480 896.000 394.040 ;
        RECT 4.400 379.080 896.000 380.480 ;
        RECT 4.000 363.480 896.000 379.080 ;
        RECT 4.000 362.080 895.600 363.480 ;
        RECT 4.000 340.360 896.000 362.080 ;
        RECT 4.400 338.960 896.000 340.360 ;
        RECT 4.000 332.200 896.000 338.960 ;
        RECT 4.000 330.800 895.600 332.200 ;
        RECT 4.000 300.240 896.000 330.800 ;
        RECT 4.400 298.840 895.600 300.240 ;
        RECT 4.000 268.960 896.000 298.840 ;
        RECT 4.000 267.560 895.600 268.960 ;
        RECT 4.000 260.120 896.000 267.560 ;
        RECT 4.400 258.720 896.000 260.120 ;
        RECT 4.000 237.000 896.000 258.720 ;
        RECT 4.000 235.600 895.600 237.000 ;
        RECT 4.000 220.680 896.000 235.600 ;
        RECT 4.400 219.280 896.000 220.680 ;
        RECT 4.000 205.720 896.000 219.280 ;
        RECT 4.000 204.320 895.600 205.720 ;
        RECT 4.000 180.560 896.000 204.320 ;
        RECT 4.400 179.160 896.000 180.560 ;
        RECT 4.000 174.440 896.000 179.160 ;
        RECT 4.000 173.040 895.600 174.440 ;
        RECT 4.000 142.480 896.000 173.040 ;
        RECT 4.000 141.080 895.600 142.480 ;
        RECT 4.000 140.440 896.000 141.080 ;
        RECT 4.400 139.040 896.000 140.440 ;
        RECT 4.000 111.200 896.000 139.040 ;
        RECT 4.000 109.800 895.600 111.200 ;
        RECT 4.000 100.320 896.000 109.800 ;
        RECT 4.400 98.920 896.000 100.320 ;
        RECT 4.000 79.240 896.000 98.920 ;
        RECT 4.000 77.840 895.600 79.240 ;
        RECT 4.000 60.200 896.000 77.840 ;
        RECT 4.400 58.800 896.000 60.200 ;
        RECT 4.000 47.960 896.000 58.800 ;
        RECT 4.000 46.560 895.600 47.960 ;
        RECT 4.000 20.760 896.000 46.560 ;
        RECT 4.400 19.360 896.000 20.760 ;
        RECT 4.000 16.680 896.000 19.360 ;
        RECT 4.000 15.280 895.600 16.680 ;
        RECT 4.000 10.715 896.000 15.280 ;
      LAYER met4 ;
        RECT 464.895 17.175 481.440 325.545 ;
        RECT 483.840 17.175 502.945 325.545 ;
  END
END user_proj_example
END LIBRARY

